�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������w������������������������������������������������������������������������������������������������������������������������������������������������������������������������������:vt�ӧN�:w��������������������������������������������������������������������������������������Ν:�p�Ç�ӧ�������������������������������������������������������������������������������������:t�ӡÇ8p�Ç9ӧN���������������������������������������������������������������������������������������ӧN�8p�FFFFFFFFFAÇ�ӧ������������������������������������������������������������������������������������s�Çdd[2-������ӧN�����������������������������������������������������������������������������������:t���Å�t���ӡÙ̂��Ý:t������������������������������������������������������������������������������������gN�:t8p�aafE�# �����N�-���t9ӧy����������������������������������������������������������������������������������ӡÇ�ȶdd����Ù�e��Ç�������������������������������������������������������������������������������������:t8p�afFE�## ������p�E��l�,8p�Ν�;����������������������������������������������������������������������������������ӡÇdddddd��������E��l��8p�Ν;���������������������������������������������������������������������������������C�8s##"�l�,9ӿ�����̋e�## �Ý:t��������������������������������������������������������������������������������Ν:t8p�̌��e� ���N�����ӡ̋e�ِXXp�Ν�������������������������������������������������������������������������������Ν:8p�̋e�ّ�Xs�������p�"�l�,,,8s�N�N�����������������������������������������������������������������������������Ν:t�p���̋e�# �Ν������t�s#### ���Ý;;����������������������������������������������������������������������������󳳧N�,,ȶ[-�t�������·22229ӧN����������������������������������������������������������������������������:t�ӧC�d[22t����Ç:w������E�ّ��p�Ý�����������������������������������������������������������������������������NΝ:t8p�̌�fFAÝ;������ @B����·22228p�N�����������������������������������������������������������������������������ӧN�8s#### ������t�V6p���W�3� g���C�2-��t����������������������������������������������������������������������������ӧN�8XXXY��Xs�����-���A�8�!]�s�R�T�q�e���:t8Y�l�d8s�N�;:w�������������������������������������������������������������������������t�ӡÇdddddd?����L��8�[�f�eU9� q�������·d[-������������������������������������������������������������������������������N�:t�p�aafE� ��N������i�S���)`s����TUʐD,�������,ȶddd8p�N�;������������������������������������������������������������������������ӳ�N�:,,,�ȶd������`�8���Q`�����8V���49������̋e�## �Ý:vw�����������������������������������������������������������������������;:t�p�Å��:w�����pi�T��Q�������X0�B�����t�s#"�l��8p�Ν;������������������������������������������������������������������������Ν:t�p���̋e� ��Ν����s8 ��Uʨ�UUUNs2� �UUU��5�`�2���·2-�̂�Çt������������������������������������������������������������������������N�8Y������Xs�����3����*@)U�UUM`#�Y�4cC*�*3':���,
�qKL g���:9�l�d[2�ӧg����������������������������������������������������������������������N�8XXY����XXp������+��r�+�ʪ��8F@�"�qL��3*@H�A�UUCP�j��$9����p�fE�ّ�XXp�N�;����������������������������������������������������������������������N�t8p��fE�## ��N�����FiX5�" s����5�8C4EdԂ)�B�-!|f�1T�k�UUJ��'�������9��l��,8p�N�;����������������������������������������������������������������������ӡÇ,,������9ӿ������V�2���kp+ae���i � ���V@@+�:�����*A�	���:t8Y��l�,8p�N����������������������������������������������������������������������Ν8p�FE�## ������鑚r�ᕸ����5�9� ��YA� � � � �f�_+Y����`V���������ddddd8p�Ν;;�������������������������������������������������������������������ӡÇȶdd[-��w����L�@�pg�����UU��ʧ4b��`AAAAAC\f)Y�dꪪ�4�\�@AfX�����:,����,8p�N�;��������������������������������������������������������������������Ν:t8p�Ù�e��l�9ӿ���Ù�x8��)`�����d�`)��P��� � � � � � �k��YF�W�9�UUNp,�0(V�#����C��fFAaÇ:t��������������������������������������������������������������������t���Å����e� ������΀W*��UUUNs2NheH���� � � � � � � �!����+  W3*����N -�����:�ȶ[29ӧg�����������������������������������������������������������������:t8p���̌��fAÝ����g3BB�\V�:���b�
����V�`A-!AAAAAAA����,�5���k*��s�R�j�����:9�l�dd8s������������������������������������������������������������������Ν:t���Å��w�����e���pe��DX*���fB�����f| � � � � � � � � � �ZBf�1T�QdUUT��,��������̋fFAaaÇ;;����������������������������������������������������������������Ν:t�p�â̌��Ý;�����9X5�H��Q]�e\�@$2��8�����f| � � � � � � � � � � � � �(�Yd��UT1S8@����:,�����,8p�N�����������������������������������������������������������������N�:8XXY����Xs������9B6r"��YΩ�iM!�UT�8�DVN)�5�� � � � � � � � � � � � � ����F*��`8eUU+s\dt9�l�?���8Y�����p�Ý;����������������������������������������������������������������:t8p�Å�t����Ι����@a��uUUUPŐ��3 � � � � � � � � � � � � � �!�+b��Ydꪥ�� ��\q�3C���Νd[-���Ӽ���������������������������������������������������������������gN�8p��# ����������I�V�YΪ�����3F6f|!i � � � � � � � � � � � � � �k��YF�V��UNr�p�i
�[�' �����:,ȶ[29ӧN�������������������������������������������������������������N�8Xs#### ��N�����I�S����ʪ�����8G`IR+c0!i � � � � � � � � � � � � � �!�+!2��YU�eNsJWʐD9BC����C���fAaÇt�����������������������������������������������������������������:t8p��̌������;����A%�T��+p,2���`i@a[�»UUT0NsH��AAAAAAAAAAAAAA|f)R4APeUUUPŁ�8��
Kg���C�������������������������������������������������������������������ӧN�8XY�����s����t,� -3�8��Җ�UU9�� �"5�
2��UUk@CK("��AAAAAAAAAAAAA�[Q����*�����TU�D a����·22-���t�ӿ������������������������������������������������������������:t�p�Å�̃�w����C��2��+�TX*����ND��-�� p�ª,UU9� +�Ns)�5� � � � � � � � � � � �`e���V��5�UUUUUPƔ��+!����N�22228s�N�����������������������������������������������������������;:t�ӡÅ���̌���;����r� Zg �*�L�UUUK �#\rKQl?�2��(p�]�UUT+Y_Ye�� � � � � � � � � �!��)e
q�k*������r�,*��X Ì�H������̌��fAÇt9ӳ����������������������������������������������������������N�222-�t����Ö �CT��Q`�����*�9 9���br�C� �TX*��̜@VN)�AAAAAAAA-!|M�0q�k*���� ��p�K,Ӆ@k���s�R�T�!����:9�l��,8p�N�;���������������������������������������������������������ӳ�·,��ȶdd������3�'$��\Җ:���9`Tʹ�8x ���:+��8��9�UT0V����S_ � � � � � � �����4@VY�eUUPŮkŠ+ ��5Hj�Ì��r��ʪ�����B�-������ȶ[29ӧN���������������������������������������������������������N�8p�##"�l�,9ӿ���t9l�+��r�Wg:���9`iB�8$�Ý���C�%�D*E|Җ
���,��4EHf`AAAAA-"�A��+ !�@Fꪪ��aV�
q�A�B�!R�Q�-�Z�US��*��H������C��̌��Çvw��������������������������������������������������������:t���Ç22-��fAaΝ����� 9X5�H�XeUUS�ҕ��8� 	2;���[-Ex8�,UU9��Zʧ43R3 � � � �� �`╓D��fNuUUT0F��Uʴ�MR�B�!B�*��*�\�e����`iJ��k�P�������fFFFAaaÇt�ӿ������������������������������������������������������w:t�p��Ù�fFFAÝ�����#4���n�ꪪ����p�,��/����#4��T��a�UU5�8CJ����AA-!�[�5�򵙐ʪ��`�*��r�,�����!B�!B�@Yf��`eUU@��8gW�������dd[28s�N���������������������������������������������������������:8p�afE�ّ�s����t�f���p�2��UUS�҄3��C��2������� 8@`,UUfB�si���HB�-!3*F�U8TfNuUUT0F`+�r�40��!B�!B�!j�AV�p��e�eUUU@)���b���:9�����Xp�Ν:t������������������������������������������������������vt�ӡÇddddd9�������qN3HWe����`�@0�A�	;�����:$��V�YΪ�����hf�k�3��
� �UUUC S4�ha\!B�!B�!B�!W
�U��
�X�����vV��!�e������ȶd8p�N��������������������������������������������������������Ν:t�ӡ���̌����;����Y�"���UU9����"�%��������g "*�TX*��k���R,���Ad��UUC�Z9e��j���!B�!B�!B�!WR�*Ҿ e����9]�2�8�x
Ka�����̋e�# �Ç:t�������������������������������������������������������N�8Xp�# �������t8XYӰ9�����9`U@)R�X�������������
�UUP�8G8��#��:���`ƼT�Ae�ePj��!B�!B�!B�!B�!WaV@S�*�`���`iJ���������ȶ[-���������������������������������������������������������ӳ�N�:8XY����Xp����3NP ���9i�YΪ���SJ��9%���������r�l�E\Ҝꪪ����Z�h
�)V�A�WB�!B�!B�!B�!B�!B��M8T�����Y[���g������̌����Çt��ӿ��������������������������������������������������t�ӧN�ddddd9ӿ���t�$�*���2�i!e��
��UT��\��$������������Qi�P$҆UUUUUC�V�W��j���!B�!B�!B�!B�!B�!B�UW8���UT��3������̌�fFAaÇt9���������������������������������������������������NΝ:t8p��̌���Ç;�����@x8!�g:�9`iM)Ϊ�9[�0(W��[����������hD*�UUUUK\���Y&�\!B�!B�!B�!B�!B�!B�!B�,�Ӗ�^-uUTҜǝ:w���:t9���l��,8p�N�:vw�������������������������������������������������N�8p�# �## ������t,���(p���,UUUP,������������Ö�J��+�:�����U�$�!B�!B�!B�!B�!B�!B�!B�!Wa�U¹^�]US��,̋e�� ���?����p��l���8p�Ν�������������������������������������������������:t���Å���̌�Ý;����C���$
2�T��UUUUT�@��g;���������	@�����a`�������h+��+�!B�!B�!B�!B�!B�!B�!B�!
�^K$�¹`��W�A�8�H�8����l9����C���fFFAÝ:t�ӿ�����������������������������������������������Ν�:8p��̋fFAaΝ������j9 P� �0UUUUUU����f���������а��"#���)Ϊ�����Z�h5�Y&�B�!B�!B�!B�!B�!B�!B�!B��f��UT+r�i
�,�ҕ�pH������p�"�l��,,8s�N�;�������������������������������������������������N�ddddd������-�%`��������	Q�*��b�N)^�/�������XIf�+sJ����  ��ʪ���V�W8�a\!B�!B�!B�!B�!B�!B�!B�PU�\� 2�����L8@AfX�����,ȶ[22t�ӳ������������������������������������������������N�,����,8s����[3NP�p��Xꪪ���T�4s�,�HT mUUNsJ�"�-Fs�������а�i�C�W�)`��� 
�Ъh͜aX���`�pY%y+�!B�!B�!B�!B�!B�!B�¬�����`ʪ������3T��9�������̋fFFAaÝ:t��������������������������������������������������:,,�ȶd����Ù��A� X*���`9S-i���L80
k�h栨@�eUT0�P  [�������e��C�W�)`����*Nq'4��4
�ak`�%hT&������b�*�^J�B�!B�!B�!B�!B�!W
�Y!
4�L-pʪ���@ʪ��L��T�Ql?����p�E�ِXXp�N�:w����������������������������������������������;:t8Y�l�d����΅��`A�J�Җ
���c^*e�4r�lЀ)�y�*F���D�UUNsJV�
�������̀�$
�\���Ϊ��cX�M9�sJ�i����]%t��ZF�������\
�9V�A\!B�!B�!B�!B�!B¸UZU¢���*��  ���g�ʈ@���`iB��`$9������̌�fAaaÝ;�����������������������������������������������:8Y��l,?����Y��+攰UUUC �L���j�5��y�y�pf�e�0UUR�+s���4?����̀�`� 0� ꪪ�b�
��\Z�
�AAJ�
�@ʠӕeUUC e�+Yd��!B�!B�!B�!B�+�0�*�X��k����Q9�Uc8#�Y4A3*���vi ��U l�������FFFAaaaÝ:vw���������������������������������������������Ν�[-������K2��W�(eUUT0T�Z�U�<��<��<��<��)��,���*��b��R�
B�����23B" $�ڪ��s�Vf �SJ�AAAA3+@� UUU-r�r�U�PWB�!B�!B�!BØU��4�L-uUUT *&����PP�B�As�q��
���4�\��f�����:,����8p�N�����������������������������������������������N�[-�̎����g �
�|Җ
���`����9�4 
y�y�y�y�y�M~V@�HT&�����YW8�R-Fs����A%�qN3HWa�UUCTV�jji]� � � � � �WEtjhPV����UUT0T�8B�$�!B�!B�!B��J���r���UUM`�Fsp��B�
(P�PpF�+%�� UUC��8x-E������̌�fAaΝ;���������������������������������������������·2-�̎���[-G$
2�iK ʪ����Q4��rVh@��<��<��<��<��<��<�
hEH��ZT l2��f�D,������Y� Zg�+p,�UUU9�2�V�y@4AAAAAA�AL�
Ш@5UUC{
�)VNa\!B�!B�+�p�`)�`����*&��8E��B�
(P�B�
As�hAQ5�UU,)_*A,�C����:t9�l�,8s����������������������������������������������ӡ�̌����t9lr@��U�a]�ꪪ���P���8eH��y�y�y�y�y�y�y�y�Њ�����UU9���8`P�,C��:t�Z�L��C*��UUT1�Z
Ъh� � � � � � � � ��ii8 UUPŮ�2�U�PWB�!B�����9h5�����Ph���((P�B�
(P�B�
(P�hPpF�9���@�2����Y�N�����:ȶd�ӿ���������������������������������������������Ç-��a�������-UUUkHYg�`<��<��<��<��<��<��<��<��<��83g�� ���]�C���4?�:g-Ex���2�UUU5�AZA�+РhW@� � � � � � � � �%tjik`�
ШNuUUC�h
ŖhR�!CT�Bi¢���UUC����0�PP�B�
(P�B�
(P�B�
(U4(8Vq���UUR���S�l�3����t9�l�,8s���������������������������������������������Νd[,Kg�Ζ��`� 0��eUUT�HYf�W0�y�y�y�y�y�y�y�y�y�y�pf�@�� UUC0$��~�Z�I�*@)S,UUSX�s�6fB�AAAAAAAAAA���S0@0* �UUK\�a\��iT��T�
���@G5�ʪ���pr3@p�)�M(P�B�
(P�B�
(P�B�
(P�B�A�#�Z��UU����$)2;���s"�l,9ӧ��������������������������������������������t�s"ٜ���Ζ�Ӕ" $�eUUP�l�J���9Y4�
y�y�y�y�y�y�y�y�y�y�y�y���d5BUUNsJ�"���p�8BC�YS,uUUC�B���� Ю�AAAAAAAAAAA�549�V*YUUPƼZ8q�ie�r�k��UUNp����DT�pESJ(P�B�
(P�B�
(P�B�
(P�B�

��D��k*��XP���?����e� ����������������������������������������������:,�X�����K0 �&�,UUC������ɦ�y�y�y�y�y�y�y�y�y�y�y�y�y�#G5D�UUCenj�B�V �� »5�UUMb�
�І`�F���] � � � � � � � � � � � �%tWB��5�h*��b��e�#�e�UUT�3%@Z��4#�

(P�B�
(P�B�
(P�B�
(P�B�
(P�B�@PpG4�����UT����B�f�����B�� �N���������������������������������������������Ν:ȶX����BJ�q@��4�����`�9S-i���gy�y�y�y�y�y�y�y�y�y�y�y�y�y�y�Y�*��UUR�4�)W4���UUT1�@a�@4AAAAAAAAAAAAAA4�PV�VUUCUUT0`����AT҅
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

��T� ,UUX2�8@@ ����[-��;����������������������������������������������̋e�l��k�ª,UUP�9S-i���Vh@��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�B*��YeL���:����QZ�aA��L+�AAAAAAAAAAAAAAAA+�SJ�2���P�������TNFq�X�((P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P(.p�a�ʉk���ҕ�T
�49��Ι�e��N���������������������������������������������C��L��Ü�0�UUU��ց� Uf�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�S�j�YP�UUUUP�h+B�+b�
�� � � � � � � � � � � � � � � � � �Ѧ��0UUUUU*%����PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

��dY�UUU, `q@�l��Ù��p�N��������������������������������������������Ν:�g	2��f��*��5 a�*�B<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��82�YeB������I�+Ѧ�� � � � � � � � � � � � � � � � � � �ѩ����UUUUU*�pAAB�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�����8�9QUU9���T�q���-�%� �N���������������������������������������������C�������l
R������0�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y��͕�G4�mUUUUP�J�B�AAAAAAAAAAAAAAAAA����@��V�BUUUUT̜�������
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

Ўa�� @UUNr�' �2�尒ِp�����������������������������������������������e�Io�3�B����b�*橯�)�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�����9kJ��UUUUMcN@�
�t � � � � � � � � � � � � � � � �%tWF���f
�V�Pk*�����Nhi�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(E8G��UUK�j����L�L尳�����������������������������������������������e�Il���
����`��s�l�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y��
ᣕr�*6UUUUUP�*f4��AAAAAAAAAAAAAAA4�8±h5�UUC �B�UUT�*&��!�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

� ����i ���23��aa����������������������������������������������C�����[�MUUUP6ZZh
���<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��0�IWYP��UUT1�+r�UU9ʄ�
�fLAAAAAAAAAAAAAA4(+b�+B�k*���eD�Y�������UUP���ӂ

(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P(*EEUUUʑ����尰�g��������������������������������������������:,�X�����`P*����l����J��y�y�y�y�y�y�y�y�y�y�y�y�y�pf�*F���AQa�UUKJV�I��@8e|��� ±T54��AAAAAAAAAAAAJ�
�A�Pʪ��*HU�R4#�4"�h�*`8eUUCPq� �(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

)�3*���]����$�[w����������������������������������������������p��b[��f��*�cX�UUP�Bj�<��<��<��<��<��<��<��<��<��<��<��<��)�Y�Y�* l2�������9D9BL��` �j��,�UUC aQ�V�A��t � � � � � � � � � � � ��
k��aPUUT��AkM�` ��y��R�4�B�UU�@������
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
p
�*���vj��� ���Xs�N���������������������������������������������:[,BKg專iSX+��-����*H�_�S�<��<��<��<��<��<��<��<��<��<�� �Uf�j
��UUCT� ��!�[w�-�%�p���9�UP� T- *� � � � � � � � � � � ��P(+c�4�B*���eD���U�<��<��<���9kJ����@TM9�p�L

(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�@F��4�D UUUT5@��e�Il,9���������������������������������������������t,ȱ	-��A�*�
�fW��*ʪ�4��VM~O<��<��<��<��<��<��<��<��<��<��0�AS�ڪ��s�P
T�q�
L��� ��UG:���Š�f4��AAAAAAAAA��MW��
�0ʪ�����,��T��y�y�y�y�Ug�� UUP�d!`aR8@PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P(8!���
�������f��2,BKfAΝ���������������������������������������������:dg,Kg專Vꡊ��
Za@��V�Q�����r�,��6pg�y�y�y�y�y�y�y�y���h�\� �YUUU,
����P� 8���Ӓp�,UT1P��^L�i��] � � � � � � � �ѩ���``V �*���ʙW4r�i���<��<��<��<��<��0�Ahj��� 9�9��
(P�B�
(P�B�
(P�B�
(P�B�
(P(8Vq����
�����U+�T�����̃���������������������������������������������Ν23�����a��C�`QE-0 �
�UUʙe����<��<��<��<��<��<��<��83ep�J�P`mUUU,
�!�3�*� ���Ù�S\j�0,2���aX��i�L+�AAAAAAA44ҽӉ4�BUUT0Z@j�83�<��<��<��<��<��<��4"�hZT�pʪ��*&��*��@PP�B�
(P�B�
(P�B�
(P�B�

��DT���`+�V����,�	-����������������������������������������������Ç23����  ��C���ER���0* �uUT0-\�
���<��<��<��<��<��<�5�R8e�i �6�������3�fp������` �T���9�UT
�2� �W@� � � � � �WEtjh2���h5�*���	�,��Uf�O<��<��<��<��<��<��<��<��0�!P��UUC +#8 ��B�
(P�B�
(P�B�
(P�@�(��4�D�����b�V�PfX-`EB�Wf��2,BKfA�����������������������������������������������:dg	-����[��+C0(��(���k��aX ���l����Y��y�y�y�y�x4"�8e���a�UUMb��I�P�#����:[-ER8E\҆UUP�
���
�AAAAJ����3��UUU�2֜IR5�<��<��<��<��<��<��<��<��<��)�ʑ������ʪ���Q4�暘(P�B�
(P�B�
(P�B�A��-d�ɬ���`+g4��4
�
ش*�f��		-��:w���������������������������������������������8s#8Il��ȪEn���F�EQEQE
�sN$ӕeUUeD�9R4#�<��<��<��)�Y�,�PZx2���b�'"�il�����t�rN	*��UUMb�V�j5ƚPAAAA+�J�l�
Š�UUU@r�Z�G5M�<��<��<��<��<��<��<��<��<��<��4"�9�*����b��,���PP�B�
(P�B�
(E*G�*!�������k��� �WElZJ����A!%�����������������������������������������������C��Kg�ERj�ZjQEQESM���Ӊ4�BUUC	�4r�k�
y�y�pf�@-iS�*����Dk�HR[;������9' �B�UUC	�+ɘ-04AA4(T�h5�UUP6TMAe�2�5�<��<��<��<��<��<��<��<��<��<��<��<��������UUP���ӂ

(P�B�
(P(8#�sY* UUT1P�c�9��i�t �%tsKB�j��� ���Xp���������������������������������������������ӡ̌�&s���j�Z��QEQEQE-`(T�h5�UT0j ²i���)��+&�ZҦ�UUUJ�sT
�9l?�����Ù�S\p������V*����� �W@T-`�
�UUP�l�J���9R5�<��<��<��<��<��<��<��<��<��<��<��<��<����W*`8eUUNr�i�2�8(P�B�A��4F���UUT0�^L�k��� � �	]�*�٪��2,BKfA�������������������������������������������������g;�2+�_UJ�b�(��(��(��(����V�� UUP�9PY�l��G-iS�UUT1`UE|���Ý�������-�!�W�(eUT0@eliT�J�l�
�����-�
ɦ�y�y�y�y�y�y�y�y�y�y�y�y�y�x4�T��!P��ʪ�  ����S�PA���� uUUC�B�$� T+�AAAZJ����a%�l,9ӿ��������������������������������������������C��L���I_UV�-1EQEQEQE�E-0 ���YUUC �L���* ,����, ��8g � 8s��������-���8E\ҜꪪEh�HV-�eUUC��j,��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�� ��*F�Z���*��Ph�aR*G05D�UUUAZ����t � � �	]�hU�P?�[w��������������������������������������������:9��$�w��uT�(��(��(��(��(��ZaA�6q�A���5�UUU9���8gU#�$�����������I��%L�UUSX�K@s����*HYf��`<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�6r�i �ʪ��ʉQ*%D ���b�+B�+`��@�AAAA
شT5@���b[2t����������������������������������������������Νdg	3���9%}T0V+b�QEQEQEQEQE���0l�
�������enq�P�r��_��������s4�C�i
�UUUUUC �L��9Y4Ã<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��)��G-iha�UUUUUP�*fLAAAA4+bЪWf��	,Kaa������������������������������������������������fp�8�Y�*�V+b�QEQEQEQEQEQE*�^��HV+�Ϊ���X@0��f����������9����X*����ʉ�@���y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�peVh
�P �UUUUMb�V�P0�
�tW@� � � � �%tVšT5@���b[w��������������������������������������������:8Y�$��rJ��i�ii�(��(��(��(��(��(��)kz9�
����Ñ�4�9����������XI�5@�UUUUT�UgO<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�� ��5KZ������0�6k�4
�AAAAAA+��-
�vj��� ��ِs���������������������������������������������C�23��!������r�-1EQEQEQEQEQEQER�H敠@����L���?����������8RrN�4�:������Hr� ��y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�N��¡UUUT�-hU �W@� � � � � � �R�-�+�T����̃����������������������������������������������:t9��$��r���V+b�QEQEQEQEQEQEQE4�@�aR����������������3J��*E\ڪ�����e��� S�<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�� ��+��Z���UUP+���(� � � � � � � �Jش*�f��tȱ	-�w��������������������������������������������:t9��$��r���V9��(��(��(��(��(��(��(��(���5�UUUT���9 p����������NP �����UUPʪ��ʙe��83�<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��83g��AP��UUPŠ�
�0 
�t �� � � � � � � �R�-
�Y����Kِs���������������������������������������������C�2,BK���*�Q��QEQEQEQEQEQEQE�E
$ UUUUCPqJ�2�������Ù�$�0��UUU-s^-Qh �\2�����U�U��y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y���p��ZT�x2���kb��@� � � � � � � � � U+bЪWf��2,BKfA�����������������������������������������������̌�%�_���*�X斘��(��(��(��(��(��(��(��H����5�UT�4�|��R[;��������fiX5Ʃ_4�����b��aQW*�@q�p���eUT0b�5�W~O<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<�
hF�@�ʀ��������J讁AAAAAAAA*��h�j���Ķ?��������������������������������������������t�s"��,B��K0$�U
�����(��(��(��(��(��(��(��(Pq �Y|+PG�UU9�)_*@@ �w��������r�"���`UUPŮ�3N��9�p��T�@P�Y�eUUT!
ɯ�)�y�y�y�y�y�y�y�y�y�y�y�y�y�y�M~W����UUUU@05i] � � � � � � � � ��lZJ����E�Il�9����������������������������������������������Ù!%�_�Y�!�-1EQEQEQEQEQEQEQE(8�U8��l��+Y�UU@��j��̶w������-�L�eniC*��0F���g0�!B��d��NZUUC �L��SL ��y�y�y�y�y�y�y�y�y�y�y�y�y�y��Y�,��*ʪ����P��AAAAAAAAAJ譋@e@�T����&p��N��������������������������������������������·dg		�:Y�g:�Tl��EQEQEQEQEQEQEQE8�T�e�1�R�4b� 2����[�3\r�'����:[
NH5J�U
����0�Uʴ�R�!B�+�PM9S �*���e��83�<��<��<��<��<��<��<��<��<��<��<��<�� ��V@�֖�^UUU�,�ʨV3t � � � � � � � � � hVšT��P?�d[w��������������������������������������������:t9��$$/�t�8�uR�B�QEQEQEQEQEQEQE�B�� �Mb�lc�lрC�3!�UT��� H�����#4��*e����b��eLӀ��W��!B�!BØU�\* �]UUP6ZZh
���y�y�y�y�y�y�y�y�y�y�y�SB*G�ʀ���Nh
��4EET0V3t � � � � � � � � �%tVšT5@���HIl,8���������������������������������������������p�E����2�T*6Zb�(��(��(��(��(��(��(��(Pq ��W͌c�3ed
�k*��`T���VL������i��V�vs�����x���%y+�!B�!B�!B�Y*�\-pʪ�ʄ�9R5�<��<��<��<��<��<��<��<��<��<��83L+ a�*&�eUUMb�T���B50�TӚT
���F��AAAAAAAAA�+b�P,��Ι��̃�����������������������������������������������dg		;�-G`�Z����(��(��(��(��(��(��(��H�k2��1�c�+ H�AΪ���U �䙡����t��C��)`����*�W*�T�p�!B�!B�!B�p�,��
�X-uUU@�i �T����<��<��<��<��<��<��<��<�� �Uf���02����TM9�p��SJ(0���Q�+�AAAAAAAAAAB�-
�vj����%�l,9ӿ��������������������������������������������Ù�А���2�T��B�(��(��(��(��(��(��(��h�AĀj�9_61�c�1�Ԋ�W�9�����U ����_���Y�VqR@a]����-r��Aʴ�MR�B�!B�!B�!B�!R�Q�-�eUU�e���
y�y�y�y�y�y�y�y�SL5@�PT@�eUU5 !Y��AB�
(3P��A��AAAAAAAAA@�VŠ�T5@��XHIl,9���������������������������������������������t9�bf�����'�U- j*���(��(��(��(��(��(��(��H�k�c�1�c�(�iRY_+XF*��iJ�� ����NP �en������3N�d���!B�!B�!B�!B�+�PM9S5�ʪ�*e\�Y��y�y�y�y�y�y�x5�\4�* ,2���@TNFq���@PP�B�
(p@eCc0W@� � � � � � � � � �R�-
�vj���"�$�d�ӿ���������������������������������������������ȱ	3L���
��ERQEQEQEQEQEQEQEQB�� �Mb�YC�1�c�1��#C+QZ�pʪ���38�s8 � P�0,�UUU-s^*��s��R�!B�!B�!B�!B�!BØU�\* �\2�����Z�@T�~y�y�y�y�y�y�l� �PT@ڪ���TMA�+&�pAAB�
(P�B��5�B��+�AAAAAAAAAA�[�S^5@��XIb[w��������������������������������������������:t9��$�2��X*���B�(��(��(��(��(��(��(��(q �b�YC�1�c�1�c8��hej+XUU9��5B!fg��fi�k��W4��Ϊ��b��aQ_��j��!B�!B�!B�!B�!B�!WR���\�\2��1P��G+�� ��y�y�y�y���H�ʹS�*��*&��#�
��
(P�B�
(p8eCF`��AAAAAAAAA
�lZ*���ȱ	-��;���������������������������������������������ȱ3BL����T�U- jQEQEQEQEQEQEQE�B�� �Nr�YC�1�c�1�c�)��Fd�UUP,�0(r�!̋�8@(�uUUC�T�8Y'0��!B�!B�!B�!B�!B�!B�p�,��
�X,*��� �+&�O<��<��<����XBʄ�UUT1�*DT��AB�
(P�B�
(P�sYT+j+�AAAAAAAAAA+��-
�vj��� ��ِs����������������������������������������������s#8HI��f�"�U-yQEQEQEQEQEQEQEP��@5SX��P�1�c�1�c�1��+  W,�ʪ�XC���pg��)`���#8VN2�5HB�!B�!B�!B�!B�!B�!B�!R�8G,*��`,�,�0�y�y���p��ZT�pʪ�� 9�8GM(P�B�
(P�B�
(P�sYS�*] � � � � � � � � �JشT��P?�d[2t����������������������������������������������Ù�BL��4�کP�@(��(��(��(��(��(��(��(�������1�c�1�c�1�c�H�� �Y:����0���,UUCX
�\�J��!B�!B�!B�!B�!B�!B�!B�!B¨*Ҿ�eUU@r�U���<����e�B��UUCPq�!�PP�B�
(P�B�
(P�B��5�B��� � � � � � � � � � �T��B�j���L�K�Xs���������������������������������������������ӡ̋4�-��iR+�R�*� QEQEQEQEQEQEQEQM4(8�T�+�1�c�1�c�1�c�1��Y4@V�1UUC*����^ʙ�,��9�p�!B�!B�!B�!B�!B�!B�!B�!B�p�iW
��Zꪪ���Z�@T���G-iS5�UUP�d�sp��B�
(P�B�
(P�B�
(P�pʡQ[� � � � � � � � � � �T��B�j����!%���N��������������������������������������������·dX������*@Z�P�@(��(��(��(��(��(��(��(�����|��1�c�1�c�1�c�1���XC沪�����k�+ �Y9�p�!B�!B�!B�!B�!B�!B�!B�!B�!B�j�d
�{-pʪ��M!kM 2���Q5 aR�P�B�
(P�B�
(P�B�
(P�C�i�eP���� � � � � � � � � � U+bЪWf��,BKaa����������������������������������������������N�2,BBK�IȀ�R�*� QEQEQEQEQEQEQEQE
$U5����c�1�c�1�c�1�c�H����sX2�����TU�3�j���!B�!B�!B�!B�!B�!B�!B�!B�!B��K,�`������eUUC �g0��M(P�B�
(P�B�
(P�B�
(P�@�i�*���� � � � � � � � � � �T��@e@�T�:�,KfA�����������������������������������������������:��f����$�j�T�(��(��(��(��(��(��(��i�AĀj��_,��c�1�c�1�c�1�cE�ieT�k�UUT*�WB�!B�!B�!B�!B�!B�!B�!B�!B�!B�!R�Q�-�����������S�(P�B�
(P�B�
(P�B�
(P�B�
8#��ʡQ[TAAAAAAAAA@Э�B�]���,�	-�;;��������������������������������������������:ȱ	3Kg��4��Ė���(��(��(��(��(��(��(��H���P�1�c�1�c�1�c�1�c�VŔs P�fC*��X��q���!B�!B�!B�!B�!B�!B�!B�!B�!B�!B¨�XוUUUP�d�Y9�4����
(P�B�
(P�B�
(P�B�
(P�B����U
�خ�AAAAAAAAA��شT5@��rı3��:w�����������������������������������������������̌�&il���8F�T 8��QEQEQEQEQEQEQEQM48�T�e�1�c�1�c�1�c�1�c�1�ellр@�����¦��J���!B�!B�!B�!B�!B�!B�!B�!B�!B�!Wa�i�5UUUB�i�2��AB�
(P�B�
(P�B�
(P�B�
(P�B�
.r3YPŠ���AAAAAAAAA@Э�B�]���8HIl,9���������������������������������������������9��$�-��'Ҫ�
(��(��(��(��(��(��(��(�AĀj��_,��c�1�c�1�c�1�c�1�c��١�pʪ����i�iT��!B�!B�!B�!B�!B�!B�!B�!B�!B�T�J���@eUUSX̕ VMNpAAB�
(P�B�
(P�B�
(P�B�
(P�B�
(P���eP����AAAAAAAAAJ譋@e@�T��		-����������������������������������������������wȱ3L������UP��
QEQEQEQEQEQEQEP��@5S����1�c�1�c�1�c�1�c�1�c6��UUUX`�(�R�B�!B�!B�!B�!B�!B�!B�!B�!B�p�&��±V ʪ��@T�.
(P�B�
(P�B�
(P�B�
(P�B�
(P�B���k*�G4��AAAAAAAAA
�lZ@�T�:$$�d����������������������������������������������N�2,BL����l�ʩT�8�HQEQEQEQEQEQEQEQE$U5����c�1�c�1�c�1�c�1�c�3��B����b��g�I�B�!B�!B�!B�!B�!B�!B�!B�!WR�����e�UUUC��j`PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B��Fk*s����� � � � � � � � � �R�-
�vj���#8Il,9ӿ��������������������������������������������Ù!&il���p
�T�8M4QEQEQEQEQEQEQE�@�� �M`�YC�1�c�1�c�1�c�1�c�1�el�B������U������!B�!B�!B�!B�!B�!B�!B�!\9�
q#*����D�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(\��YT�M�� � � � � � � � � � �T��B�j����Il,9���������������������������������������������9��$�-����U*��P(��(��(��(��(��(��(��(�����|��1�c�1�c�1�c�1�c�1�c��e���*�T@pʪ�Z�WJ�s
�B�!B�!B�!B�!B�!B�!B�+�d�Y�
�2�UUUUT1�9�AB�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(\��YT�@AAAAAAAAAA�[�ʁf��X��̃�:w�����������������������������������������������E�H�w�[8T�ka@��(��(��(��(��(��(��(��H����1�c�1�c�1�c�1�c�1�c9�Id*�BU������eUT0`**��+�!B�!B�!B�!B�!B�!B�+�p�`)�`�������4�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
-d U*��� � � � � � � � � �R�-
�vj���B�Ķ���������������������������������������������t8s"�$�-����SU5�2�QEQEQEQEQEQEQESM
$UW͌c�1�c�1�c�1�c�1�c�1��$�R�8f͕�G*�L���k�L��i�+�!B�!B�!B�!B�!B�!B���NT�x��*��b�*��+r����9��(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�Z�k��	�@AAAAAAAAAA��AΨj����Il,9���������������������������������������������C�!&i����
 �P�a^�LQEQEQEQEQEQEQESM
$U5�ec�1�c�1�c�1�c�1�c�1��5�B�iSf͕Y\4�T 8eUUkŠӀҨ+�!B�!B�!B�!B�!B�+�PU�\+��������T
�i� ��PƜ��
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B嬄
��恠 � � � � � � � � � ��¥R�5@��p��ِs�����������������������������������������������̌� r����
 �SX�
�(��(��(��(��(��(��(��(�����|��1�c�1�c�1�c�1�c�1�c�K!T1�9f͚a�Y\4�i
�2�����i�Up�!B�!B�!B�!B�!j��4�L-uUUR��g,��fFhD*储cNjr�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P���*�	�@AAAAAAAAAA+�0T��P?�$$�d�ӿ��������������������������������������������N�2,BL������ �S��p��(��(��(��(��(��(��(��H�k�c�1�c�1�c�1�c�1�c�1�el�B�i@ٳf͛6l�2�5B�UU,9�$�!B�!B�!B�!B�+�PU�\+�`����`UE\��`�;�' ��CsS�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B����T�@AAAAAAAAAA+�0T5@���BKaa�����������������������������������������������̌�h�;�25�1T�+B�
(��(��(��(��(��(��(��i�����|��1�c�1�c�1�c�1�c�1�c[��CC�6lٳf͛6l��j
����Z�{
ŖhR�!B�!B�!B�p�Hi�A�UUT�, qKL���2+�[��4�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
-dU-��AAAAAAAAAJ��J�Y��̌�%���N��������������������������������������������·g	�'�F��*��hk�QEQEQEQEQEQEQEP��@5SX!�P�1�c�1�c�1�c�1�c�1�c�K!U4� lٳf͛6lٳeVj���* l2����0��T��!B�!B�!
�\*��*�\�e�eUUK�+橮9BL��Ü������P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8"�BR��AAAAAAAAA���TR�5@��r�$����������������������������������������������t8s#8H�;�25�n����QEQEQEQEQEQEQESM
$U5����c�1�c�1�c�1�c�1�c�3��B�cHr͛6lٳf͛6i�ʑ�h�- l2����ʹ�W��B�!B�!B�s
�Yf���k�UUS���!�p
� -����`�����M(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B����T!T�AAAAAAAAAA+��J�Y���,Kِp���������������������������������������������ӡ̌� r���8D+pʆ+C0(��(��(��(��(��(��(��(�����|��1�c�1�c�1�c�1�c�1�c�K!T1�9f͛6lٳf͛6l��YY4r�T�pʪ�׊�W*ӘWB�!B��Ti_
��XUUT1Us�C�$/��ҰW�C��P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8#��
� �AAAAAAAAAJ��A�+�T��		-�;;���������������������������������������������ӡ̋4w�d
�U+C0(��(��(��(��(��(��(��(�������1�c�1�c�1�c�1�c�1�c�(Y
�P�U�6lٳf͛6lٳf�0����*�@�UUPƼT�9V�A\!B�+�0� ���`eUUSJV����j-����9J�eC,�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B��@2� � � � � � � � � � �ј
�@�T��,K8Xs���������������������������������������������C�-��@�!���������QEQEQEQEQEQEQEQB�� �Mb�lc�1�c�1�c�1�c�1�c�1��%�����f͛6lٳf͛6lٳf͛+���ʀ�����i�iT�p�+��d�i_
�2�UUU+�UʐD9K���t�C*�"�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�� �T!T�AAAAAAAAAA+�0*�٪�Ä���Ý���������������������������������������������C���8H�s�U4�-3MQEQEQEQEQEQEQE(8�T�+��1�c�1�c�1�c�1�c�1�c�(Y
��!�6lٳf͛6lٳf͛6lٳeVW@��T!�*������ATd
�X,*��Xenq��2���Ӕ9�MA�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
�@2LAAAAAAAAA�3R�j����!%������������������������������������������������C���8I��Ф�
�Q �MQEQEQEQEQEQEQE4� �@5P�|��1�c�1�c�1�c�1�c�1�c�hY
��9f͛6lٳf͛6lٳf͛6l٦+� ������\�eL+�r���eUU9��*�9BB����NR�s��,�M(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�� ����� � � � � � � � � �WF`*9�+�T�:$$�d����������������������������������������������ӡ̋�8I���k��2�ZQEQEQEQEQEQEQE(8�T1_,��c�1�c�1�c�1�c�1�c�3��B�cHr͛6lٳf͛6lٳf͛6lٳf�i�ʑ�9kJ�UUT1k����`,��0(rB�?����9J�eC�*�P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
��@2LAAAAAAAAA�3PeJ����Fp��Xs���������������������������������������������N�23��p����̩UR�i^�X4�EQEQEQEQEQEQM4(8�T�e�1�c�1�c�1�c�1�c�1�c�q@��UM!�6lٳf͛6lٳf͛6lٳf͛6l��#T��ZZ uUUUUU, `p�!�g����Ӕ9�J��
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�� T!T�AAAAAAAAAA+��J�Y��Ö!%�����������������������������������������������·[3���C��#�p�*�@����H���4�EQEQEQEQEQE(8�T�+��1�c�1�c�1�c�1�c�1�c�8�Id*���
�ٳf͛6lٳf͛6lٳf͛6lٳf͛*��h�- 8eUUUR�ҕ�I�w�������*�P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8#�U �U0AAAAAAAAAMM9��TҜ ��,�,KfAΝ;��������������������������������������������t�s#8I����AW�s�aX�Ni^��(��(��(��(��(��(�����|��1�c�1�c�1�c�1�c�1�c�K!T1P��f͛6lٳf͛6lٳf͛6lٳf͛6lٲ�+����3^���WeL��T�p�����f�
�@p���
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P����
�� � � � � � � � � �)Tʥn�e�Il,9���������������������������������������������9l�f��C�� +傪� ±�sKH�E�(��(��(��(��(��hPq ��W͌c�1�c�1�c�1�c�1�c�1�P$�SHr͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6We�06����C5MqX������� S�"�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P��`:���* � � � � � � � � ��`ӆT��P��9b[w��������������������������������������������:8Y�$)3C���S�W��UT0�3ez-1M4QEQEQEQEP��@5SX!�P�1�c�1�c�1�c�1�c�1�c�K!T1P�U�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٲ�h�UTҜ0 �3������� ��P�@p�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�q��P@TAAAAAAAAAC\
��U"��t8HIl�9ӿ��������������������������������������������Ù!!I��3� ���� ±�l��(��(��(��(��H�k���1�c�1�c�1�c�1�c�1�c8�Id*����6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l٦aU����X-������ $�U �H((P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B��3*���� � � � � � � � �	]L
�+ڥvC?��3��̃����������������������������������������������:t8Ybf�&h���5�UUUB �q&��
i��(��(��(��P���|��1�c�1�c�1�c�1�c�1�c�K!U4� lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6T�,UM!�-��������	9�TJ�PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
�3*� �� � � � � � � �%t��ӌ*5�J��,�����$�9������������������������������������������������E�HRf��Ü����*��@��p)��(��(��(�AĀj��_61�c�1�c�1�c�1�c�1�c�s@��Ui@ٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6i�����NH�����: KC�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�A�**��^M4AAAAAAA����f �V���9�SJp�p ���		-�:w��������������������������������������������t8s"�$)3C�Ü�J���@
�UU@a���(��(��(Pq ���(c�1�c�1�c�1�c�1�c�1��"�Ui@ٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6i��QU�������� 2�T�� ��B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8#@TUB��PAAAAAA�+�*���+	���s�enT�P��fp�ِs����������������������������������������������s"�$)3C�Μ��r�VN3PTC*��@�3 @��(��(��AP���|��1�c�1�c�1�c�1�c�1�c�hfUSHr͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳL*�@TUC%`�������Q�,TJ�PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
�**��^@� � � � � � ���05�T*���8?�rı-�������������������������������������������������f�&i���fq��D���ʑ�4�D�UUP�*�� ��QE*��UW͌c�1�c�1�c�1�c�1�c�1��fUCC�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6h�ET�8���������&�`�
�T҅
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P��QU5���AAAAAJ讍4��ią`2����]�2������̃����������������������������������������������:9��$���Ζg2�Q9� �s�3�q���k*����3 Ai�h���UC�c�1�c�1�c�1�c�1�c�1�f��T���f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�
��P�X;�������p��T�� ��B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8#@fUMb�4�AAAAA+������h5�UUUU,�t9��3��:w���������������������������������������������ӡ̌�!H/�t p�uR�s\�r��Ug�*&����Š��� ��4� �
�T�+�1�c�1�c�1�c�1�c�1�c�s@C2����f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�U�Ъ	+������2�U*%H((P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B��@ZMb�4�AAAA����B��8°k*���WeTV�UJ�ᖣ��B���Xs���������������������������������������������ӡ̌�!H/�t�8g:�Q4 �r�˗.jr�4���ʪ�k��!�L*��U5��ec�1�c�1�c�1�c�1�c�1��̪�4� lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛4«4ET0V������)8ev�TJ�PP�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
�**��Th � � �	]���+�Z��UUS��4�
�D8�R�ᖯ�9b[2���������������������������������������������dg	
@���s��@p�.\�r�˚����*&�����QZc+CYT�e�1�c�1�c�1�c�1�c�1�c�s@C2��C�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛*�@TUP$�������Rp��T�����B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8#�TUMb�4�AAA��4�G4�
�BUUR��9K"�
 �R�8e��,BKfA�����������������������������������������������:����΀PʥD��˗.\�r�ˌ����UUMb�i�9P���_,��c�1�c�1�c�1�c�1�c�3��PƐ��6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͚9QU��������3MP-T�����B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�

aQU5���AAJ����� ���UUU���8$)2;�-2�9�,2���		-��:w��������������������������������������������t�p��He�:��:�Q8�\�r�˗.\�r��p��*!����T�e�1�c�1�c�1�c�1�c�1�c�s@C2��C�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͚aU�Ъs�e`�������Ҥ���(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�s
��b�4�AACM

��B�P�UUS���`
r �Y����i�0ʕ��-_����Xs���������������������������������������������,�3L��B�T�U*&�e˗.\�r�˗.\�E�9�#*! eUUUCYe��1�c�1�c�1�c�1�c�1�c9�!�Ui@ٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l��hUN2�w������iR�J��

(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�@��P�`W@�WF����!Z��2��� Y[�g ��A��-0�s�X0��Yb[2t������������������������������������������������fE��;�
MPʥD��r�˗.\�r�˗.\��8G0�eD�UUUT*9�l1�c�1�c�1�c�1�c�1�c�hfUCC�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛*�G-
��2�w������iR�J��

(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�C�9�EU
�4�J��KH�aX�MeUUXP
p��̱�Ζ�C9�+����e�b[w��������������������������������������������:t8Y�bf���I�X*���e˗.\�r�˗.\�r�˄Q�#@r0*���9Z��[c�1�c�1�c�1�c�1�c�s@C2��C�*�f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l��Ъs�%`��������HU3'0((P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B���TUSXӁ��^@��������9%��w�Ζ�C�`p�W��	-��;���������������������������������������������B̌�!!�iR,J��2�˗.\�r�˗.\�r�˗.3�sFT���d��+a�c�1�c�1�c�1�c�1�c9�!�Ui@ٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�Ė�T	+�����f� -T9�AB�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(¢��9P�������UE�p�!�����a�+��������̃����������������������������������������������N���BB��
�d�r�˗.\�r�˗.\�r�˗.N�9���@UUP*ae��1�c�1�c�1�c�1�c�s@C2��C�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6q%ET0V�������*@Z�s��
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(P��QUUUUT�4�np�^ �G��KL!����e�bgt�����������������������������������������������s"�HH_��IȋR�h�\�r�˗.\�r�˗.\�r�˗.\"�ӘZ�Q5�UT0 �0��ح�1�c�1�c�1�c�1�c�ʪi@ٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6i�Vq%ET�J���������#J����iB�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
.Z�����s�TU�D38��:U �s�Wg�΅�!%������������������������������������������������p��bX���'",L�jr�˗.\�r�˗.\�r�˗.\�r��(�i�5����p��sF,���1�c�1�c�1�c�1�怆eT1�9f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٲ�8����%c��������UP��B�
(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
8"�UUU���8$[�����a�,2���,BKfAΝ��������������������������������������������Ν[,BB��BN`����\�r�˗.\�r�˗.\�r�˗.\�r��s
�UUU�Ej43el1�c�1�c�1�c�1�g43*��9f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳgTUC%`��������iU@s�(P�B�
(P�B�
(P�B�
(P�B�
(P�B�
(��5�UUPƔ8A�	���:Za2�vp��e�Il,9���������������������������������������������:t,�X������"�T\�r�˗.\�r�˗.\�r�˗.\�r�˜ӑ�
�����QZ���(�1�c�1�c�1�c�s@C2���U�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳfʬ�J�����������,N�U� PP�B�
(P�B�
(P�B�
(P�B�
(P�B�

��Uf�ӕUUTg��������*X0�X��������������������������������������������������N�������q@�P4"�˗.\�r�˗.\�r�˗.\�r�˗.\f�UUUUB0**���(�c�1�c�1�c�1��̪�4� lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6Uf�����IX;��������UP��P�B�
(P�B�
(P�B�
(P�B�
(P�B���4"� @����P
T�6r������t��Ω`q�?��Il�9�����������������������������������������������в�bX�����(���2�˗.\�r�˗.\�r�˗.\�r�˗��h�ʪ�-pʪ���k+Q��Q��1�c�1�c�1�怆eT0B�Sf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf����J���������SJ�S
(P�B�
(P�B�
(P�B�
(P�B�
*�9��*!Ϊ��X�rL�#�����KL!�T�@�r�$��������������������������������������������������fE�b���(��jr�˗.\�r�˗.\�r�˗.\�r�˗.\f�̪�{
�U������U���(�c�1�c�1�c�ʨ5dٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6i�Vh
��`$�������I�4���pE
(P�B�
(P�B�
(P�B�
(P�B�A����@�UUUSX��lw����:Za2�8Y�΅�!%������������������������������������������������в�bdw�[8�Z�@r3B.K�.\�r�˗.\�r�˗.\�r�˗.\f�̪�*e�U�(V�eUU�9_42�9��1�c�1�c�ʨcPVM�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͚9QU9���w��������R�@q�B�
(P�B�
(P�B�
(P�B�
(8G�*!����(O����Ö�C��g�fp�ِp���������������������������������������������t8Y�bX�����UFsK�.\�r�˗.\�r�˗.\�r�˗.\�q� T1S*��*�V��X#��UT��|eH�c�1�c�1��̪��PVM�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳfʬ�P�IX;������9�*�P��

(P�B�
(P�B�
(P�B�
(�2��2������������:Za�T�3���Il�9�����������������������������������������������p�ٜ$��-�J��sK�.\�r�˗.\�r�˗.\�r�˗.\�q�#2���i�`(V�UUNp�W��VMHc�1�c�3��PƠ��6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf�0��QU��������3��U3�(P�B�
(P�B�
(P�B�
(8G0�eD�UUU��,�Uq������t��eC����s9b[t���������������������������������������������:,�X�����UFsK�.\�r�˗.\�r�˗.\�r�˗.\�q�#2�Z�L�L0`���5�UU���Q�9��1�c�hfUC�Tٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l٠**��2�w������s�UJ��pE
(P�B�
(P�B�
(P(
ed* �UUT�3%k+Q��0C5�S��;�����Ra�5�Ô��9b[w��������������������������������������������·2,BK��4����ir�˗.\�r�˗.\�r�˗.\�r�˗.3DfUC2�0`��d�MAh,*�����eH�c�1�g43*��AY6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6h�EU8����������SU5���
(P�B�
(P�B�

���r�UUP�9dXVFf��uP��;������*X����,KfA����������������������������������������������N���L���`P��McNp��.\�r�˗.\�r�˗.\�r�˗.\�q�#2���i�0`��Z�r���UT#8�%H�c�1��̪�5dٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6i�VhB�c����������5SX��P�B�
(P�B�
(P(
V@B�*&����V�эH��A|T�֪�g����t��Ψ`0��Ù�Kaa�����������������������������������������������C��!%��� (UJ���8E˗.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`���,��M9h5�ʪ�s�r�h�ɩc�s@C2���͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf��*��IX;������9�*j���jaB�
(P�B�
(P(.p�3��B�UUU5�8�"�V�`AC_"����;�����Ra�5������b[;���������������������������������������������e��$����� �SXӜ"�˗.\�r�˗.\�r�˗.\�r�˗.\f�̪�*`4��0`���,�Y8�,����UT�,�+4EH�c�ʨcPVM�a�f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�KB���������3���k#S
(P�B�
(P(8#S��!`8eUUC���F�jF`AH����H��H�j�9�,�����:Za�T�?�9bX�̃����������������������������������������������N�-��Kg�f��*�Ɯ�.\�r�˗.\�r�˗.\�r�˗.\�r�4FeT0TU�0`��Id�0`��Yf���eUU9� 
���sNi�9�!�Uj
ɳL6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf�l�J��`$���������ESX��P�B�
(P(
�#@iʈ@���cX� ����AAB�5�R+Z�q������t�A2��Ô��9b[2t����������������������������������������������ӧB�fp����Y���i�r�˗.\�r�˗.\�r�˗.\�r�˗.3DfUC0`��0`�d��0`�d�8�,ӕ0��UT�,����l�FeT���lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6UgTUNp$���������ESX�hP�B�
*�pC+%���5�UU�k+Q����5�� � �ZF���T1������t��Ω�g����Xs���������������������������������������������t8Yl�[;�k�b�cPp��.\�r�˗.\�r�˗.\�r�˗.\�q�#2�**�0`��d�0`���Y'e�p����9dp	
沨cPVM�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳfʬ�J������������*�L(P�B�A���p*����f���S0 �� � � ��ZF���T0V������i�3�R�,���p��Xs���������������������������������������������N����%�����T1�8A�r�˗.\�r�˗.\�r�˗.\�r�ˌ��P�L�L0`��0`��0`�J�U�ӕ0��UT�3!#PƠ�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6q%ET0V�������k�"�`"�(U4��������UUT�3!QT�YA�� � � � ��k��Z�C%`�����Ζ�C�b�,���p��Xs���������������������������������������������t�Yl�[;�
�T1�8A�r�˗.\�r�˗.\�r�˗.\�r�ˌ��P�L�L0`��0`��0`���,��4�L-uUUUT1�5M�6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳfʬ�J�����������3��H�8As�hFUUSX#�@VN)�AAAAAH� �UJ������-0�s�k����rı-����������������������������������������������C����%����A[�T1�8E˗.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`��0`��,��,���`4��@k������*�f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�U���s�%`�������a�*�朩 0!`8eUUC �k+�k6fp� � � � �!i���*�J�������9%|�T�3���p�ِs������������������������������������������������E�8I�?�8D+pʆY�.\�r�˗.\�r�˗.\�r�˗.\�r��h�ʨb�U�0`��0`��0`���Y%�h
��� e�����BYeHٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6l�P�IX;������  ��R�TD ����Y#�fAAAAAAHB�
�Np$������䀧:��e�g���������������������������������������������������ӡe��$�w�+uP�@p�)r�˗.\�r�˗.\�r�˗.\�r�˗�3*��i�0`��0`��0`��$�Ld!A¹^�]UUT1S
�f͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6Uf��*�J��������n��:���V�����)���HAAAAAA-!(*UN2������NH
s�k����Yb[w���������������������������������������������B�fp�8�p ��UY��˗.\�r�˗.\�r�˗.\�r�˗.\f�̪�*`4��0`��0`��0`��,��*�B�5�E{-pʪ�����ɳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛4r���%`�������MpUUUU9� 
�Y8�`AAAAAAA��HB�
�C%`������$9�5�����9b[;��������������������������������������������Ν:[,BK��R+ꡂUe˗.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`��0`��0`��0`�K$� 4#XW,��UUT�2�h�d�͚a�f͛6lٳf͛6lٳf͛6lٳf͛6i�Vh
��c�������Ä�a�j���`�e|��("���-!AAAAAAAHB�
�Np$������䀧:�8r���Ķvw���������������������������������������������-��K��W�P��"�˗.\�r�˗.\�r�˗.\�r�˗.\f�̪��S�0`��0`��0`��0`��$����hF��#*��`6Tʹ����6i��lٳf͛6lٳf͛6lٳf͛6lٳL6h
���q�������Ö��`
2��UUk��
�[�AAAAAAAA-!(*U@S�������T�?�9��-��:w���������������������������������������������[3����Ζ�WUJ��R�˗.\�r�˗.\�r�˗.\�r�˗.3D��*`4��0`��0`��0`��0`��*�B� ��UUC��Z�G+&͛6lٳf͛6lٳf͛6lٳf͛6l�U����e`�����Ι� AȀR�,*��cX�e|�͙�_ � � � � � � � � ��ZBPT�9!�����9 )Ω�g�K��Xs���������������������������������������������t8Yl�	,C��U�*�B�p�.\�r�˗.\�r�˗.\�r�˗.\���Ui�0`��0`��0`��0`��0`�
U�ʪ��`6ZZh�d�͛6lٳf͛6lٳf͛6lٳf͛6Uf����J����������(eUUC��
��3�-"�-!AAAAAAAA��qeJ�9e���������2��r�����XYӿ���������������������������������������������вٜ$��:W��T!�.\�r�˗.\�r�˗.\�r�˗.\�q�#2���i�0`��0`��0`��0`��0`�V�r�UUUUe����j�Y�f͛6lٳf͛6lٳf͛6l٦Y�**����w����9���	�����s�@IeS\!i�� � � � � � � � � ����q
�8
W��������2��r���Ķvw��������������������������������������������t�вٜ$����2�*G �r�˗.\�r�˗.\�r�˗.\�r�ˌ��P�L�L0`��0`��0`��0`��0`��0�X*����*%�4sT�͛6lٳf͛6lٳf͛6lٳL6h
��`$��������CT!�a�UUU�fAAAAAAAAAAB�-!H�Nr�9!�����9 (eM`0�;�:X���Ý���������������������������������������������p��b�t�YΪTd"�.\�r�˗.\�r�˗.\�r�˗.\�q�#2���i�0`��0`��0`��0`��0Y%�q�b�U9��d��UU@�Q5�j�Y�f͛6lٳf͛6lٳf͛6hB��q������9b *��J�������Ae � � � � � � � � � � �ZB8�ʜ�)������XC*X���X��̃����������������������������������������������B�fp��?�rK,�U*%d"�.\�r�˗.\�r�˗.\�r�˗.\�q�#2���i�0`��0`��0`��0`��0`�N0�X*�40*3!�UP�l�MA����6lٳf͛6lٳf͛6l�U����e`����s#4�C��)`����UT
�HAAAAAAAAAAAB�5Ƥq
��S�������T0r���,BKaaΝ;��������������������������������������������:t8Yl��t�XeR�VB)r�˗.\�r�˗.\�r�˗.\�r�˗��CEZ`��0`��0`��0`��0`��,��+
�� ���R9� W3!�UT�P�Vlٳf͛6lٳf͛6i�����8�����Ι� AȀ�Wj���-r��0�X*��P� � � � � � � � � � � ��!�B�`0������Ӓ���ag��,K�Xs���������������������������������������������t�Yl�f�����s���K�.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`��0`��0`��0`��0Y'V,P�YC[�Y �*��b�5 a�T��a�f͛6lٳf͚aU���s�%`�����H8e|҆UUT1��P�d
宪�Y�AAAAAAAAAAAH���*�\������9 )Ω`g���l�9ӿ��������������������������������������������ӧB�fp����X8�*��p�.\�r�˗.\�r�˗.\�r�˗.\���UT�i�0`��0`��0`��0`��0`���T��P�1����� �UUP�D���R6i��i�͛6lٳfʬ��P�IX;��g,���2�UUPŁ^¢�J���@5T
�(AAAAAAAAAAAB�Ԏ!U+��������3���p��Xs���������������������������������������������t�Yl�f���Μ��U*'0�.\�r�˗.\�r�˗.\�r�˗.\�q�#2�*�0`��0`��0`��0`��0`��W,Nr�YC�1�敓Dq�k*��b�5�rH��0��6lٳfʬ��P�IX;���#4��T���ʪ�0FsP�T��5@i^�P+,�AAAAAAAAAAAHCR8�T�������9 )Ω�g����XY���������������������������������������������:,�g		����TNa�.\�r�˗.\�r�˗.\�r�˗.\�r�4FeT1S*�0`��0`��0`��0`��0`�d�a\�UJ�ec�1����De�s���� 搲�@�ʬٳf͛6i�Vh
���q����� �UUC�r�*�T��!
�,�P�VlAAAAAAAAAAAB�Ԏ 2�_�����r@S�SX,���Il�9�����������������������������������������������p��bf���)��TN`˗.\�r�˗.\�r�˗.\�r�˗.\"���R�*eZ`��0`��0`��0`��0`��,��+�
�9_,��c�0�1��R@��*���T%@Yg T��6lٳL*�@TUNp$���V ��f��UUP���j,�¸B�!W id*�VYB � � � � � � � � � � �!�Z�W���������2��e�g�L�%���N���������������������������������������������N�2,LА��Ӕ�U*&�e˗.\�r�˗.\�r�˗.\�r�˗.\f�̪�*eZ`��0`��0`��0`��0`��,��+�
��e"�c�1�c9�H	��s���b�4��pʑ�f͛*�@TUC%`���r�8@a�,UUZ�TU�iT�!B�!
�,�T�(� � � � � � � � � � � ���
�R�U ��������T0Y��e�b[w��������������������������������������������Ν-� s4��9NΪTN`˗.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`��0`��0`��0`��0Y'W,C2��1�c�1�g4�%|#�ʪ�5�pʑ�fʬ�P�IX;� 9X5Ʃ_4�����x�����!B�!
�*ª#\ � � � � � � � � � � � �
�*�� ?����Μ�2��Y���3����������������������������������������������������e���3B��@�ΪTM ˗.\�r�˗.\�r�˗.\�r�˗.\���UTʴ��0`��0`��0`��0`��0Y'W,Nr�YC�1�c�1�c9�H	��k*��`,�,�#eH*S�+p�pT�(UUC�^¢�U�PWB�!B�!
�*¨c�*B � � � � � � � � � � �!��P�|������KK 0�;�g	-�;;���������������������������������������������dX��&_�j*E���4.\�r�˗.\�r�˗.\�r�˗.\�r�4FeT1S*�0`��0`��0`��0`��0`�d�gX*���1�c�1�c�3�sJ���G5�UT0*�4�j ڪW�!�,$�C�V�2�������40��!B�!B�p�J���r�k�AAAAAAAAAAA�XeNr�U ��������T0Y���,BKaaΝ���������������������������������������������C���9�e��� -T ir�˗.\�r�˗.\�r�˗.\�r�˗�3*���V�0`��0`��0`��0`��0`��a\�U9�e"�c�1�c�1��S�Y@k+��UUP�9h- mU@����p��HWj���-p**�ZU�B�!B�!B�aU
�HAAAAAAAAAAAA8�VT�������9 )Ω�g����Xs���������������������������������������������t�Y�bf��_�Yi��P���r�˗.\�r�˗.\�r�˗.\�r��h�ʨb�U�0`��0`��0`��0`��0`��W,P�YC�1�c�1�c�1�� 5��ʪ�����!�3JUUPƼZ@
U��WB�!B�!B�!\8�B�ʐ� � � � � � � � � � � �q@�U+p�������C*k%���rı-���������������������������������������������ΝdX��i��tqJ�T�5���\�r�˗.\�r�˗.\�r�˗.\���U-p��0`��0`��0`��0`��0`��a\�U9��ec�1�c�1�c�1�� 5���k*��������{
�8,��B�!B�!B�!BÌ�*�\��AAAAAAAAAAA8�VT�� �����-2�R�8e��g	-��;;���������������������������������������������:dX��i��V�����Ӏ\�r�˗.\�r�˗.\�r�˗.3DfUC@4��0`��0`��0`��0`��0Y'W,P�YC��1�c�1�c�1�c9��he|�f�eUUUUUUXp��d���!B�!B�!B�+�hU�\ � � � � � � � � � � � �!��n�����[��UP���b[;���������������������������������������������N��&h/�����T *'#9�a�r�˗.\�r�˗.\�r�ˌ��P�L�L0`��0`��0`��0`��0`��0�X*����1�c�1�c�1�c�1�g���A�UUUUUPŮ�3NU�Pj��!B�!B�!B�!B�q��T*+" � � � � � � � � � � �![0ʆ+p�������r��,���9bX�̃����������������������������������������������B�e��-����EUP��si�.\�r�˗.\�r�˗.\�q�#2���i�0`��0`��0`��0`��0`��q���W�(c�1�c�1�c�1�c�1���42�As�������j R��¸B�!B�!B�!B�!BaU+YY5� � � � � � � � � � � �2�P�n�����C���i5���	����ِs�N���������������������������������������������C���4[���S�Wj����a�8˗.\�r�˗.\�r�ˌ��P�L�L0`��0`��0`��0`��0`��3�,P�YC�1�c�1�c�1�c�1�c9��hej
�0�UUUK\�aQW��j��!B�!B�!B�!B�!\8�B�V�� � � � � � � � � � � � �R��n����̋Qi����)�W�q�w��,BKaa����������������������������������������������ӡfE��-��T�UUP� �0��˗.\�r�˗.\�q�#2���i�0`��0`��0`��0`��0`���S�!�P�1�c�1�c�1�c�1�c�3�l���V�YUUXp��g0��!B�!B�!B�!B�!B��5T*+&�AAAAAAAAAAAA)_�V�����9bY�4��,��Ù�KaaΝ��������������������������������������������ΝdX��r��t�%����� 
ɡR�˗.\�r�˗.\f�̪�*eZU�0`��0`��0`��0`��0`�N0�X*�e�1�c�1�c�1�c�1�c�1�c8���q����3PJ���!B�!B�!B�!B�!B�d��U+YYAAAAAAAAAAAA(C9�J�"�����')�5Jܮ�uT�B!���3���Ý���������������������������������������������B�e��-��@@US��UUP� �dЂ)r�˗.\�r�ˌ��P�L�L0`��0`��0`��0`��0`���q�r�T0C,��c�1�c�1�c�1�c�1�c8�`暑��A�T*�PWB�!B�!B�!B�!B�!B�%�2�Z�ɮAAAAAAAAAAA@�U9ΪV�/���t�rN	�vs���|�����Ķd?���������������������������������������������[,L�9l��� �T̜A�@eUT1�* ��r�˗.\�r��h�ʨb�U�0`��0`��0`��0`��0`���8¹`�����1�c�1�c�1�c�1�c�1�f`��PU-s�,��!B�!B�!B�!B�!B�!\*�SUB9��AAAAAAAAAAAC9�M!�2���t� 
�W*��UUT�+����3��̃����������������������������������������������·[	3KQl���8�v�kA��De�UUfJ�+&�\�r�˗.\f�̪�*eZ`��0`��0`��0`��0`��,���P���1�c�1�c�1�c�1�c�1�c�i��B����B�!B�!B�!B�!B�!B�Y*a�B9���AAAAAAAAAAAA)T�:��_��V ��+�UUUT5@��rı3��:w��������������������������������������������:t�Y�H)-����]��aT��jEd�A�9�UT̄,���K�.\�q� T0TU��`��0`��0`��0`��0`��I��S���P�1�c�1�c�1�c�1�c�1�c�4b�UU���!B�!B�!B�!B�!B�!WS����� � � � � � � � � � � ����0
��L�Q�8�,UUUT1e�g�e�Il,9���������������������������������������������t�p�"�2;�t�8 Z��V���sJɢ8�2k*��jR58E.\�q� T1S*�0`��0`��0`��0`��0`�d�a\�UV�R�1�c�1�c�1�c�1�c�1�c8��UJ�h�!B�!B�!B�!B�!B�!B��*a�B9����AAAAAAAAAAA3S��0
��3� ��U�)������Q* mU9ʸB��,BKaag���������������������������������������������г �8����8�T#
�ec�H�� �fNuUT1�5R58E.\f�̪�*eZ`��0`��0`��0`��0`��,��+�
�9Z��c�1�c�1�c�1�c�1�c�1�S�UJ�h�!B�!B�!B�!B�!B�!B��
�*�sC5�i � � � � � � � � � � ��E*��T05�_�:$�5�����UUC �L��9�5 mT1WC���b[;;��������������������������������������������Ç2,@�Il���8�T#
�ec�qMH����UUMc2jU����@T1S*�0`��0`��0`��0`��0`�d�a\�U9���c�1�c�1�c�1�c�1�c�1�S�UJ�h�!B�!B�!B�!B�!B�!B��
�*�sF5�i � � � � � � � � � � ���B1T��C/��rN( �UUCf�5M����S���!��s9b[t���������������������������������������������t�p�"������iUNr�YC�1�c5#�s2UUTMA�VN`B�eP�L�L0`��0`��0`��0`��0`���q�r�T�+Q��c�1�c�1�c�1�c�1�c�1�0T���B�!B�!B�!B�!B�!B�!\,��2�d��HAAAAAAAAAAA��(
s���(e�:g,�!ȀR�X*���AkM���y� Z*����9�$����������������������������������������������:t9�l��%���84��W�(c�1�c+b�9�(T�UUMb�T  UC�`��0`��0`��0`��0`��,��+�
��Z��c�1�c�1�c�1�c�1�c�1�ӘUJ�h�!B�!B�!B�!B�!B�!B��
�*�A���AAAAAAAAAAAB��)�� ����hB�T��j���ʙe�2�83�<��9�P�|�;�X����Ν���������������������������������������������N���@�Il���k�*�F��8��1�c��ԍ�r���UUUUZ i�0`��0`��0`��0`��0`�N0�X*�+Q�c�1�c�1�c�1�c�1�c�1��F
�R�J�B�!B�!B�!B�!B�!B�@TT��� � � � � � � � � � � ��E*��U�P��K`s�p0Xꪪʄ�Y�`<��<��9Ъs�s���9��-��������������������������������������������������̋8Rg;�-��J��\��1�c�1�c+cR9�)Z�02�����@0`��0`��0`��0`��0`��I��P�|Ԇ1�c�1�c�1�c�1�c�1�c�h�U- 4�!B�!B�!B�!B�!B�!B@TPŐhf�AAAAAAAAAAA��(
s��S�gÖ� A�*攰���eD�9R5��y�y�r�U+�)���8Il,9���������������������������������������������t��尐8Rg;�-��J�k2��1�c�1�c8��+X�����@,��0`��0`��0`��0`��0`���q�r�T�+Q��c�1�c�1�c�1�c�1�c�fi�uT#���!B�!B�!B�!B�!B�!s�k��A�����AAAAAAAAAAB�"����`p�S8I�k�C4��UT1�e�2�80
y�y�y�j��ʆ+�)��s9bg2w���������������������������������������������:,ȱ��9��l�R��e�1�c�1�c�1�R�42�F����U��&$��0`��0`��0`��0`��$�
傩�V�c�1�c�1�c�1�c�1�c�1�gт�T#�i\!B�!B�!B�!B�!B�!B�Ak��A�����AAAAAAAAAAB�� ���S�p�3HWj���*PYg l��<��<��<��<�-
�9_9N�Ù�9�Yӿ���������������������������������������������p� �8Rg�2�T�kAec�1�c�1�c[Q�����eUUK�i�q�,�0`��0`��0`��0`��$�
储b��1�c�1�c�1�c�1�c�1�c8��V�T� ��!B�!B�!B�!B�!B�!U\��K ��|ZB � � � � � � � � � � ���UR�*f�2����ZZh�p����<��<��<��<�*a�J���t�X�̃����������������������������������������������p�E�)3����MT�8��1�c�1�c�1�c�,�C+�Tk*��k�aQ�QVLI�0`��0`��0`��0`�d�gX*�+Q��c�1�c�1�c�1�c�1�c�1�1Z�P�HB�!B�!B�!B�!B�!B�!T@eP	3� � � � � � � � � � � �!� uUUUU�2�pʬ��<��<��<��<��<��@�*�*�)��s8I�,8y���������������������������������������������ӧB�e�),N�����U5� ��c�1�c�1�c�1���42�Y�UT��0�Uʴ�%�`��0`��0`��0`��0q�r�T�+Q��c�1�c�1�c�1�c�1�c�2�4b�UB8!B�!B�!B�!B�!B�!B�P�]TL�� � � � � � � � � � � �R�ʪ����p���d� )�y�y�y�y�y省QU9��B��3�&s �����������������������������������������������C�-� p��;��MT1�!�c�1�c�1�c�1���,�C8�UUR�+�W*�4�&0`��0`��0`��0`���+�
���lc�1�c�1�c�1�c�1�c�1�����P�U�p�!B�!B�!B�!B�!B�!B�8��U��AAAAAAAAAAA���������Q-i��#_�S�<��<��<��<��<��<�-�J��w�t�X��Ý���������������������������������������������B�e���'����kAR�1�c�1�c�1�c�VƤhaPeUUR� ¹W*�0`��0`��0`��0`�
傩�V�c�1�c�1�c�1�c�1�c�1�gъ֪�pB�!B�!B�!B�!B�!B�!
�+��h��� � � � � � � � � � �f(g�����r�U�U�<��<��<��<��<��<��<�-�J��w�t�g2w���������������������������������������������B�e���!����H��
��1�c�1�c�1�c�1��Z�eUUU,
��5���Y&0`��0`��0`���q�r�T1Z��c�1�c�1�c�1�c�1�c�1�SF+Z��iB�!B�!B�!B�!B�!B�*��Z�9�3 � � � � � � � � ��ik�T��AΪ��*&���@� S�<��<��<��<��<��<��<��@�T1_C��r��d����������������������������������������������t8Y�b
K���V�8W+#�1�c�1�c�1�c�3� ꪪ���YX��iVK$��0`��0`��0`�
傩�V�c�1�c�1�c�1�c�1�c�1�g�J�h�p�!B�!B�!B�!B�!B�!B�5���#0 � � � � � � � � � �`═*3*���l�������)�y�y�y�y�y�y�y�r�T�*�w��X��Ý���������������������������������������������·[,LФ��U"�9�B��1�c�1�c�1�c�1�c5 UP��UPŁd`�J�`��0`��0`��8� �U5��lc�1�c�1�c�1�c�1�c�1��ªUKAV��!B�!B�!B�!B�!B�!C�j]T4F`AAAAAAAAA5�5#C+�Tk*���9�4���<��<��<��<��<��<��<��<��@�U*�)��s9bg2w���������������������������������������������:,ȱ3B�����V�9¢�V��1�c�1�c�1�c�s@B�UB �+�ʪ�b��X8�I�0`��0`��gX*�+Q��c�1�c�1�c�1�c�1�c�3�s
�U- 4�!B�!B�!B�!B�!B�!B�PZ�8fAAAAAAAA5�E*F�� �UUUP6ZҸpg�y�y�y�y�y�y�y�y�y� Z*��!���9bg2;���������������������������������������������N���B��?�9^
�Ϊ��c�1�c�1�c�1�c� �eU
����-�UT�*�VJ��&0`��0`��8¹`��F�1�c�1�c�1�c�1�c�1�c�)�R�Z iB�!B�!B�!B�!B�!B�9����M`� � � � � � � �����s
�
� 2����S9 
y�y�y�y�y�y�y�y�y�y��ʜ�\!�Ù�L�aΝ;���������������������������������������������:,�,C�Μ��s�*+%l1�c�1�c�1�c�1�el�P�hZB�`�%hZ*��`�@
q�0`��0`��,��+�
�9Z��c�1�c�1�c�1�c�1�c�1�SF*�T� ��!B�!B�!B�!B�!B�!sAk���!�AAAAAAAH���42�V�YUUUUC�g�y�y�y�y�y�y�y�y�y�j�0ʥ|�;�:g,L�A�����������������������������������������������p��I�X���9%|2�9Z��[c�1�c�1�c�1�c� uP�hW�M4�����A����,9�,���&0`��0`�d�a\�U9��lc�1�c�1�c�1�c�1�c�1�S�h�R�Z iB�!B�!B�!B�!B�!B�9���U�C0 � � � � � � �`eH	8��9�UU-r���l���<��<��<��<��<��<��<��<��<��<�T
����w�t�X��Ý;���������������������������������������������C��4��:rJ�eR��1[c�1�c�1�c�1�c�x2��ЯB�h���P2��r����,9�,���&0`��0Y'W,Nr��1�c�1�c�1�c�1�c�1�c+cF*�PŠ���!B�!B�!B�!B�!B�!a�,M`� � � � � � ��3���k�*��b�+�S
��Z�b�k��<��<��<��<��<��<��<��<��<��+%L2�9W9N�Ι�L�A�����������������������������������������������p��bf�!��NIW9�J�s
�c�1�c�1�c�1�c�hfUMb�+Т�)��Za@����0eUP�ZAe�eY0`��@`��$�8��T1Z��c�1�c�1�c�1�c�1�c�1���R�Z iB�!B�!B�!B�!B�!B�9���U�C0 � � � � � �`����p������b�*�d�XG�ks_�y�y�y�y�y�y�y�y�y�yY* ʥ|�;�:g,L�ag��������������������������������������������t�s#8Ib�t�s�P�Ts1�c�1�c�1�c�1�f��P�hW�EQE4�M-`(Tr����¦i�,�4�Y%�`��a\�UV�c�1�c�1�c�1�c�1�c�1�"�S�*����!B�!B�!B�!B�!B�!C�i�SX3 � � � �!��VM�A����c^*f��I�B��Z�l�����<��<��<��<��<��<��<��<��<���S�b�r���3�&s ����������������������������������������������8s#8Il?�V ÝT#�1[c�1�c�1�c�1�c� �eT�+B�QEQE�KL(Ěr����5�i�,�4�`��a\�UV�R�1�c�1�c�1�c�1�c�1�c8��UJ�h�!B�!B�!B�!B�!B�!B�&��U9��fAAAB��Ә�A����`W��Uʴ���+ɧ,C��<��<��<��<��<��<��<��<��<��<�� eNr�r���3�&s �������������������������������������������������FrĶ�@0�U,�F+a�c�1�c�1�c�1�c5 ̪�+B�
(��(��(���iӉ
�BUUk�LӖY�`��a\�UV�c�1�c�1�c�1�c�1�c�1�gъ�U- 4��!B�!B�!B�!B�!B�!s9`�s��� � � ��ZBfH���G5�UUX`+ �Y5HB�!�i�yT1kM0��<��<��<��<��<��<��<��<��<���P*�|��:g,L�A����������������������������������������������t9�l�3����PŐh�l1�c�1�c�1�c�1�g4,�P�hW�EQEQEQE-0�g a�UP�T�8q�*�3�,Mb��1�c�1�c�1�c�1�c�1�a�0T���B�!B�!B�!B�!B�!B�!a�,Nr��AAC_�#�,��UUR�5��i�iT�!B�5M9�*�-i�y�y�y�y�y�y�y�y�y�yY* ʆ*�)��s8I�,8y���������������������������������������������t�s"�I�/�t! �YT���1�c�1�c�1�c�1�怆eT1Z���(��(��(��)k�V��UU-s^*e|�f$�B��UV�c�1�c�1�c�1�c�1�c�1�g�J�h�p�!B�!B�!B�!B�!B�!CTӄb��V�0 � � �`ԎaT�Q����k�a\��g0��!B�+ɧ�Pŭ4��<��<��<��<��<��<��<��<��<��+%@S���!���9bg2;;���������������������������������������������Å��8��8�CA���1�c�1�c�1�c�1��fUMb�-!M4QEQEQEQE+��8 �UUK\
��B����`2�b��1�c�1�c�1�c�1�c�1�a�1U*�- 4�!B�!B�!B�!B�!B�!B�\וNr��A���42�U@:���� �j,���!B�!R�kʡ�Zi��y�y�y�y�y�y�y�y�y�VJ�2�W9N�Ι�8Xs���������������������������������������������:t9�l�3���3��U,�C8��1�c�1�c�1�c�j@!�UV�zQEQEQEQEQE-`�F�0����k�eL+���UC�Ԇ1�c�1�c�1�c�1�c�1�c�)�R��iB�!B�!B�!B�!B�!B�5J��*��j� ��8�H�YdUUT1��N��5HB�!B�!
�W5�Pŭ4��<��<��<��<��<��<��<��<��<��+%L2�W9N�Ι�L�A����������������������������������������������t8Yl�3����X*�A��P�1�c�1�c�1�c�1�ԀC2�k�^�QEQEQEQEQE�����UUC�eUV�R�1�c�1�c�1�c�1�c�1�c8��UJ��8!B�!B�!B�!B�!B�!B��_5�T
�i�C0qJ��ʪ���^¢�q�¸B�!B�!B®kʡ�Zi��y�y�y�y�y�y�y�y�y�VJ�T1_C��r��d�����������������������������������������������d[,L�����,Lɡ���1�c�1�c�1�c�1��̪�+B�
(��(��(��(��(��(���k���P������j5!�c�1�c�1�c�1�c�1�c�Fh�k9�KAV��!B�!B�!B�!B�!B�!B��וP�����he|#���UT1`U��Ye�W��B�!B�!B��W5�Pŭ4��<��<��<��<��<��<��<��<��<��+%@S���!��s9bgvw��������������������������������������������·-�%���8e���43R�1�c�1�c�1�c�3�B�b�+Т�(��(��(��(��(��(���``Tk*���s��R�1�c�1�c�1�c�1�c�1�c���U- 4�!B�!B�!B�!B�!B�!B��yU9�9Z��8��5�UUkŠӀҨ5HB�!B�!B�!�U�yT1kM0��<��<��<��<��<��<��<��<��<���S�W�S���r��d���������������������������������������������Νd[,K�� p�S2��01�c�1�c�1�c�1�ԀC2��HQEQEQEQEQEQEQE(3����UUUC�c�1�c�1�c�1�c�1�c�1�g4ъ֪��WB�!B�!B�!B�!B�!B�5J��*�cX����k��+�r�*��B�!B�!B�!B�U�yT1�6y�y�y�y�y�y�y�y�y�y�d�uCs���霱3������������������������������������������������p��bX���T�U3 I�c�1�c�1�c�1�c�ʩ�V��Zb�(��(��(��(��(��(��(��`@`Tk*��*Y��c�1�c�1�c�1�c�1�c�(��j�h�!B�!B�!B�!B�!B�!B���UUUUCX
�)VMR�!B�!B�!B�+�\UMAU�y�y�y�y�y�y�y�y�y�yY*S���!��s8I�,9ӧ���������������������������������������������Y�l�,B���X*��$Ԇ1�c�1�c�1�c�1�怀:�b�+Т�(��(��(��(��(��(��(��h�A�!Z�YUUM`�9��(�1�c�1�c�1�c�1�c�1�ӘV�T#���!B�!B�!B�!B�!B�!
��Z*�������N��+�!B�!B�!B�!B�\וC��y�y�y�y�y�y�y�y�y�y�d�R�r���-�&s ���������������������������������������������:ȶX�!� �,@p$Ԃ(�1�c�1�c�1�c�3�B�b�-!EQEQEQEQEQEQEQEQE�
ШMeUT0 �0Ԏ(�1�c�1�c�1�c�1�c�sM�j�G�!B�!B�!B�!B�!B�!B�hA`����k�aQW8��WB�!B�!B�!B�!
�W �SPT�<��<��<��<��<��<��<��<��<��<�� eC����$�����������������������������������������������t���E��$/� �Z����1�c�1�c�1�c�1�����hZB�(��(��(��(��(��(��(��(��)i�`�!X�UUP�d*
ɩ��1�c�1�c�1�c�1�c�9�kUB9V��!B�!B�!B�!B�!B�+�PU��׃*��1`U��Yf��%p�!B�!B�!B�!B�5@PU5Vy�y�y�y�y�y�y�y�y�y�d�Nr�r���3�&s ���������������������������������������������:ȶX�!�Rr"�U��R�1�c�1�c�1�c�3��SX�
�(��(��(��(��(��(��(��(��(��)i�±����c2�B�jC�1�c�1�c�1�c�1�g0�g:�G�!B�!B�!B�!B�!B�5K$5�����c^*f�!E�j��!B�!B�!B�!B�!P�j��AR<��<��<��<��<��<��<��<��<��<�T�J��w�t�[;���������������������������������������������C������)9]���I�c�1�c�1�c�1�c�ʨb�+Т�(��(��(��(��(��(��(��(��(���*����8�DVMH�c�1�c�1�c�1�c[1U*����!B�!B�!B�!B�!Wa��AV ʪ����ʹV���!B�!B�!B�!B�!B���T1�*G�y�y�y�y�y�y�y�y�y�VJ�eC���9��3�:w��������������������������������������������Νd[,K/�r"�U5��Q�c�1�c�1�c�1�g43*��ЯB�(��(��(��(��(��(��(��(��(��i��f8eUUUf@���R�1�c�1�c�1�c�VƌUJ�h�!B�!B�!B�!B�!
�\*��*�PZꪪ�� � S@W��B�!B�!B�!B�!B�!B���U5Vy�y�y�y�y�y�y�y�y�y�d�*s����9�$�d�����������������������������������������������dg,BL��9Ȋ�T��c�1�c�1�c�1�c�ʨb�-!EQEQEQEQEQEQEQEQEQER�U����d+�"�jEl1�c�1�c�1�c�qM�j�h�!B�!B�!B�!B�!�Y !�-�2���W��U�B�!B�!B�!B�!B�!B��j��*G�y�y�y�y�y�y�y�y�y�VJ�U+�(���I��9����������������������������������������������:,�dw�f� -T�Hc�1�c�1�c�1�c�hY
�9Z�i�(��(��(��(��(��(��(��(��(��(�@*�D���UC�q��Q�c�1�c�1�c�qM�j�h�p�!B�!B�!B�!B�s
��r�,*����ep�!B�!B�!B�!B�!B�!W R���4�H��<��<��<��<��<��<��<��<��<���PT1W9N�Ù�KfAΝ�����������������������������������������������e���/��8�Z��V���1�c�1�c�1�c�3� ꡊЯB�(��(��(��(��(��(��(��(��(��(��q�j���9�!P
��s�@���ьc�1�c�1�c��R��iB�!B�!B�!B�­*�Q^�\2������d��!B�!B�!B�!B�!B�!P�j����y�y�y�y�y�y�y�y�y�yY* ʜ�|!�Ù�Kaa�������������������������������������������������fr�$����8�Z�`���(�1�c�1�c�1�c�3� ꡊЯB�(��(��(��(��(��(��(��(��(��(��q�
����i�9�!P ꪪkp��#�1�c�1�c�1����U�4�!B�!B�!B�!�h,�3^���]�Q�5�PŠ�+�!B�!B�!B�!B�!B�!B���2���� S�<��<��<��<��<��<��<��<��<���PU*�)����Il�9���������������������������������������������·23�!&_��q@�T�C61�c�1�c�1�c�1��U5�д�QEQEQEQEQEQEQEQEQEQKH� �Mc��p�sJ� uUU9�9_YR9�c�1�c�1��1U*��HB�!B�!B�!
��4 )�`��*��cJW�S�p��`�#�d!B�!B�!B�!B�!B�!B��j�P��<��<��<��<��<��<��<��<��<��+%L2�W9N�Ö�KfA�����������������������������������������������Å��L�#��4��kF�����1�c�1�c�1�c�ʩ�V�z�EQEQEQEQEQEQEQEQEQE(8�SX��S�.\"�ҲZ�QUT��|e�V��1�c�1�f�UJ�G�!B�!B�!B¨8ʸT��eUU,
�
p���g� ��d!B�!B�!B�!B�!B�!B��R�+���<��<��<��<��<��<��<��<��<�T
���B��-��̃�;���������������������������������������������N�2-������5�T��c2q�T�h�1�c�1�c�1�g3*��ЯB�(��(��(��(��(��(��(��(��(��(��q�j�����r�˄S�sFTBUU5�9_YeQ�c�1�c�4`�U-ZB�!B�!B��d�(��^���9]��$��9��r�*�h8��\!B�!B�!B�!B�!B�!B�uT��
y�y�y�y�y�y�y�y�y�yY* ʆ*�)��s8Il�9���������������������������������������������·-�������
���G+�YEl1�c�1�c�1�g43!�9�д�QEQEQEQEQEQEQEQEQEQKH�Mc��r�˗й�8G0��k*�������Q��1�c�qM�j�h�!B�!B�!�*�
ʰXUUP�Y_*A�	��HT#�ep�!B�!B�!B�!B�!B�!W B�U4�p��<��<��<��<��<��<��<��<��<���PU*�w��[2t����������������������������������������������:,�f����&�4��� �dԆ1�c�1�c�1�P̪�+B�
(��(��(��(��(��(��(��(��(��(���Āj� jr�˗.\�r�8F��`�UUP�+YT�YGc�1�g4ъ֪��WB�!B�+�PU�\*+�k�UUSX��Äfs��+ b��2�B�!B�!B�!B�!B�!B�+�4�
��+���<��<��<��<��<��<��<��<��<�T�uR����a&s �g���������������������������������������������p��H���	-2�V�v�����4EH�c�1�c�1��%���
�(��(��(��(��(��(��(��(��(��(��ZG@� �.\�r�˗.\��8F��eD�UUP�+YZ����ac�qM*UK@!B�!B�W��Q�-�UUR�4��9 p��r�*���+�!B�!B�!B�!B�!B�!B�aU4�p��<��<��<��<��<��<��<��<��<���S�b����a%� ���������������������������������������������:,�	��C�!�����b�+�YGc�1�c�1��D�C�i
(��(��(��(��(��(��(��(��(��(���Āj� jr�˗.\�r�˗.p�4�D�UUSX�`)�,��1�c8���R�HB�!B�s
�YaX�e�UUKJW�S\r�Ý�Õ�%U�ZWB�!B�!B�!B�!B�!B�p*�eR�+���<��<��<��<��<��<��<��<��<�*a�W����8I��9���������������������������������������������·-�&i�g;��Kg()Ϊ�k��r�jEl1�c�1�c8�Id*��hZB�h��(��(��(��(��(��(��(��(��(����*� !�˗.\�r�˗.\�r�8F�ӕYUU�P
s���3�h�R��iB�!\9�ZU ��*��`i@S�U"�g���`�Y 4��!B�!B�!B�!B�!B�!
�U�T����<��<��<��<��<��<��<��<��<���J�U+s��t�X�̃�;���������������������������������������������C��4)	w���NI�+�v��8�����1�c�1�P$�C�^�QEQEQEQEQEQEQEQEQEQKH� �B ��˗.\�r�˗.\�r��Ug�*&���
��9���g4aU�
+�!CT�K,Ӗ�����`i0(r@�G��+ J�Y 4��!B�!B�!B�!B�!B�!
�U�T�����<��<��<��<��<��<��<��<��<���UJ����-�&s �g���������������������������������������������p�Fs4��9����Pj��`��� ���(c�1�c�K!T�+B�
(��(��(��(��(��(��(��(��(��(����*� !�˗.\�r�˗.\�r�˗.2�8�AQ��� ъ��0�U@2�j��+���b��UU4�|�����:��Y 4��!B�!B�!B�!B�!B�!aU*f��y�y�y�y�y�y�y�y�k�U�uU+s��t�g2w���������������������������������������������C��B�����dY�C���UU5�9T�YEl1�c�qMd*�+B�QEQEQEQEQEQEQEQEQEQE
0T N\�r�˗.\�r�˗.\�r��Ug�*!�UT
��+��Z�L!E�Y%ZU¢�������S 3����)ƪ�@+�!B�!B�!B�!B�!B�!B�����3T�y�y�y�y�y�y�y�y��
ɣ�@UP�rC�Ù�KfA����������������������������������������������t�p��H Z���s9b:[+��S�UT�@!Y5"��1���d*�+B�
(��(��(��(��(��(��(��(��(��(����*�  ˗.\�r�˗.\�r�˗.\�r�*F�!e{5�UP��UR�-X������83�rLг����,�5T� i\!B�!B�!B�!B�!B�!B�ZR�j�y�y�y�y�y�y�y�x6r�T 8eUR�V�Ù�KfAΝ;�����������������������������������������������e� Z����r��?�3J�r"�,UC��42�sF1�elh�!T1Z���(��(��(��(��(��(��(��(��(��(Pq�j� 2�˗.\�r�˗.\�r�˗.\�s�jr�8�A�UUUUUZ�2��s�e|������t�8�R�
�B�!B�!B�!B�!B�!B�ZZR�W<��<��<��<��<��<��<��٠-iha�UP,�?�尒�Xs����������������������������������������������:,�X��PR[;��3J�V� !�*g:��b�+�YC�Vƈ�Mb�+Т�(��(��(��(��(��(��(��(��(��)ia�@�r�˗.\�r�˗.\�r�˗.\�s�jr�h�A���������*�� ����t�8j�d ��B�!B�!B�!B�!B�!B�ihUJ�Y<��<��<��<��<��<��<�B*F�Z��k��UT�,� ���3��̃�;���������������������������������������������ӡ̌�h���Ak����9l/:[9@�iUUSX*Jɩg	,�P�hW�EQEQEQEQEQEQEQEQEQEP�� �B ��˗.\�r�˗.\�r�˗.\�r�˗.MNV@���
������X��8$e����r��9�J���!B�!B�!B�!B�!B�!BihUJ�Y<��<��<��<��<��<��)��P0�6����)_*ER	;���!%� ���������������������������������������������·23�����Ф5�$�,N��P8	9'��j���8�$��� ���s��^�QEQEQEQEQEQEQEQEQEQKH�@p��˗.\�r�˗.\�r�˗.\�r�˗.\�E59Y4E@fC*�����4�|�5�`$?����Ӕ�UJ�Yf�B�!B�!B�!B�!B�!B�ZZR�j�S�<��<��<��<��<�6j���*��b�*�" _��l$�-��;���������������������������������������������ӧC��L�����V ��9KL�2�)�Á��T�
��� ����Y���HQEQEQEQEQEQEQEQEQEQE(8�5P�59r�˗.\�r�˗.\�r�˗.\�r�˗.\��4#�h� UUUT�*����w����:Y�0ʥ{MR�!B�!B�!B�!B�!B�!\*�Ъ�� ��y�y�y�y�pf�@��02���L8�$�;��K4$������������������������������������������������C��BK�p V��x+hB s��2 ㌩�UU5� ��uT1Z���(��(��(��(��(��(��(��(��(��)ia�@�r�˗.\�r�˗.\�r�˗.\�r�˗.\����� ���b���9&i������: 8g:�^�ST�!B�!B�!B�!B�!B�!W ihUJ�� S�<��<��<��<�U�֖�^���vi3�VB���f���Xs����������������������������������������������:t8Y�$$��+!�ҩ����S8s�Ι���@�UUUP�hW�EQEQEQEQEQEQEQEQEQEP�� �BDhE˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.NiY  @���a�5�(H�����@�ΪW��5HB�!B�!B�!B�!B�!B�p�K@eR�r ��<��<��<�
hEp��AQa�UT�+sT��!��Ù��ib[w������������������������������������������������!&_�p9X9%`����$�! �$���ii����ڪ����hW�EQEQEQEQEQEQEQEQEQER�8�5P�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˚�\"�#�i�uU9���@@ ������t p�uP+�!B�!B�!B�!B�!B�!Be�U*' O<��<��<�
k�T5B�UT�4�\�B��w��t���s ���������������������������������������������������E���/�t�9J�rB�H�,B��W��,N�����p�!`����
�(��(��(��(��(��(��(��(��(��(��ZG�#B.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗80���[� ������� ��@0��!B�!B�!B�!B�!B�!
��T�*��<��<��<�6r�T 8eUUU@)�Q���:$�!&s �����������������������������������������������vt9�l$�3���B�e�fL Y���� AaΙ�P*�ʪ�+��EQEQEQEQEQEQEQEQEQE��0�T 4F�\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗50"����eH w������@�U �R�B�!B�!B�!B�!B�!B�+�Y*j�Q9 
y�y�U�2�T��eUU+��S������%����l,9ӿ���������������������������������������������C���L��?���Q�9%`"��@� 	,�2��t��9'��a�UR�8��k�(��(��(��(��(��(��(��(��(��ZG@��#B.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗8d*�n������: 5NuS^*�B�!B�!B�!B�!B�!B�Y*a�J�� S�<�
peH��ZT@ڪ���8��B�;���� 
BL�A����������������������������������������������Νd[	����3��(D9'$#eR	�+�.d3C�9T���,0c�P�B��-1EQEQEQEQEQEQEQEQEP�� �BDhE˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r� ��ES�9'�����:Z�����sT�!B�!B�!B�!B�!B�!C����D��S_��0�UUP�XC5B6r�!���:d  �9b[t�������������������������������������������������e�X���r� ����A�+�f�,J�X-��Y��i( P-T
�P0 SMQEQEQEQEQEQEQEQE��0T �r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\���s�%`�������9R,@0�!B�!B�!B�!B�!B�!B�%MUʹU����j
�2���4�\�@Af[;�����p8 �-@p�9�s����������������������������������������������Ù��9�dw���)+�^ ���f�� r�~t�r��
�
���JІ`QEQEQEQEQEQEQEQE��0�T 4F�\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗50����+�����:*E��U�R�!B�!B�!B�!B�!B�!
�T�*�D���\� uUUK�"��/���̌�h � �9�g-��;���������������������������������������������Ν2-������r�),�� [9KL�,J�^ 峿Ö���I����Z �ez-`QEQEQEQEQEQEQEQE
0T4F�K�.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r� ��EP�IX;�������9R,@2�W��!B�!B�!B�!B�!B�!
�T�U`8`ʪ�X �$✓4,����L��pfY�P$�-�:t����������������������������������������������:�ȱ3KPRe��Ä���X�%�r��2����	;��a!�UP� V8���(��(��(��(��(��(��(��)i`�@r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\��+ T0V�������"�T׊�^HB�!B�!B�!B�!B�!B�p�KB������vi9K���Ö�KQfY�e� )3BK# �N�����������������������������������������������a�̌� pj	-���Ö�e��
@�A��AT�_�� �QΪ�b�4�y3 @��(��(��(��(��(��(��)ia�@h��r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.ja�+ U8��������΁ʑ`�k�|�$!B�!B�!B�!B�!B�!B���UUUT���38����fij e�f 
@�%���,8s�������������������������������������������������p�#8HR  �����8RV2��9  ��8s��9N)_,UMb�V��qT�QEQEQEQEQEQE(8�5P�4"�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�s�V@"�c��������*E���r���!B�!B�!B�!B�!B�!\*�W-uUUU9�(
p��l����L�8 �9K0  ��Г9l�,8s����������������������������������������������w�:,ȱ3B�f 3L����Yb I�V3.t�Y�g���9�UB ��Ni^�LQEQEQEQEQEQE(8�5P4"�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�s�V@"��q���������3NDX*��_+�B�!B�!B�!B�!B�!C�U�Nkʪ��� ��Ze������L�8 �9K2� ��Г9l�8s�N����������������������������������������������:t8Y�l$�
@�f 3Ka����3NS�ˇ ��;��f �JUT 4�j����(��(��(��(��(����*��e˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r� ��EP�IX;������$��r���!B�!B�!B�!B�!BØU�*5�ʁf��UJ�g ������Z�3��,�0 R		,KfFAaÝ�������������������������������������������������̋e������,�PHY���8r� !|,��� w�rĬR����-hl�ERQEQEQEQEQE(8�5P��r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\#C�V@ eC%`�������Wj��W��B�!B�!B�!B�!B�!\*����00e@�$�+�`�vi�9L������r�Ij,�S�� ��X�̌�Ý:vw�����������������������������������������������Å���9j g)f����󥰐�В�9 r�$����H� ��UT - a�
QEQEQEQEQKH� �@pЋ�.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r��)Y �����w������I�+�S^+�B�!B�!B�!B�!B�PM9h5�ʪ �X5�`C*�H,�����:�f�3��,�0 R3BK�l�,8s�g����������������������������������������������t���Ù��8R ,�2� [���̎R��3NS�Y��-�f��4�:����a@��(��(��(��(���*��!�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r��Y ��V������	8@Z�`i�R�!B�!B�!B�!B�%����X*���	+R+� �w���e� Y�e�f -AH�	,KfFAaÝ:vw�����������������������������������������������t�p�E�9bf��P �9K2�w��峒W�9l),��T�L);�:g+��UUT�J�F`QEQEQESM�@`@� ��.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˄hp
�U���������	8Ev�X��B�!B�!B�!B�!
��*�
��Z�UCp�[·;���9�b,�3��,�HR	,L�s# ��Ν;������������������������������������������������N�d[3�&hRZ��fY�������"��R���U  �-�%�_�p��*EnWj���@l�E�
i��(��(��(��
� 2�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�s�V@"�����������N`�X����!B�!B�!B�!
��8ʸW �*���*�$�����s ���9K2� Z��9�X��e� ��Ν;:w�����������������������������������������������;Ν9��l�	��fr�`4������I��)X5�AfY����?�@ ��eL2��@H�QEQEQE+�*� !�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r��Y ��V������3�P-T�50�!B�!B�!B�!\9�Ziʙ��eUS�+�H��N����[3@��Y�`���BK9l�,,8s�N�������������������������������������������������C�2-���9j g)f 	;��� �� F�HBH��$䖠��s��p-UU*NW�0
(��(��(�zP�59r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\#C�V@"�`$�������[8 Z�`j
�B�!B�!B�!CT�j9`UUiJ��-2�dw���г8 Y��)f -@p8HI��dd8s�gs�������������������������������������������������:t8p�"�b
KQfY�e�Rg���fifZe�rNI�	,NI�+��9�Zg"+r�UT1h+Cf���EQEQJ� j�8jr�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�s�V@"�����������g U,9�!B�!B�!B��V@P�U��2����'� s/���E�R 9NR̳,�PX���Aa�Çt����������������������������������������������������N�,�g,BL�� ,�2� f����� 9j9NHB��@ _���6p�`eUSX*8�ش�LQEQE+�*� `˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r����ES�	+������� �Xr���!B�!B�!a�U� �e����vi9!!���Ö���9NR̳ ��X��fAaaÝ;;��������������������������������������������������t�p���ٜ$$Z�2��,�PI�����l�9NIfr@��/�-�����S��S�UT4�j(��(�zP�p��.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�F�+ T0V������3� -T�
�0�!B�!B�+�0�*�L����XC8f�!�����[	-E��r�e� � p���dd8s�g��������������������������������������������������ӧC�d[3���Ij e�f�����K� V +����`�3B�Ä����`���JІ�QE+�*�  ˄h\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�ˌ��EP�IX������3�J�XAT�!B�!B¨*�NZ02��҄3T ����:�f�3��,�0j��%���d9ӧs���������������������������������������������������w:8p�"�b
@�fY� ���Ι�`��  ��P �$��"��0�UU5�@sKH���@`@� ��.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗Y*!����������� Ҫ�U!B�!B��YaX��eUT�4�)�*�j-����t,� g)fY�`�3BK9l�,8s�Ν����������������������������������������������������Ν,ȶg,L�9j g)f 	2��[ ��� ��3NI�3L��+���󥳔
&�UU ±T(-3\V���@��r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\���	+��������SU, �B�!B�*�
ʰX*��b��
L���Ι� ��,�0j
@�hIb[-��t��������������������������������������������������������:,,ȶX���Ij g)f�!g� &\�RW��8r�䕃����	9'��ڪ�b�+@5�A�B ��˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r� ��EP�IX;�������k���k�AT�!B�­*�\-uUU,
���f����[	
K3��,�0j��K9l�d8s�N�����������������������������������������������������N�9�l�X��fY��4���N��I�9!&s4! ���䖠���p�p�!`���`� UB e˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r� ��ES�	+�������qSU-p�U!B�AV�p�׃*��8V���p���·-�����9K2� ��ВĶ[22�s������������������������������������������������������:t�p�fE�9b-E�fr�` �#���,���r�
�W�4$䕃?�t� �I�9�UC*� �.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗8d*�J��������F������AB�*�����UPƔ�� � -����t9l� �)�Y� �g-�̂Ç�ӿ�����������������������������������������������������N�,ȶg	3B�� ,�R�),B���XHR �+$$��V)_�UUU A�.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˜�C%`������� (T�K\+�AWR�,��+�`UU9�(
p�L�����:g�S��,�  �f���fAaaÇ:w�������������������������������������������������������ӡÙ�e��
@��Y� �p���8p��r@��������A�iUUT \�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.p
�U��������̍qSU-p�Y$9�W
�{-uUT1�U@I���9����r�H r���f -AH$�3�̌�Ý:vw������������������������������������������������������t�ӡÅ����H) e�f 	-�����Q�9%x+�Rw��ȳ�UUUT�9��˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�p�V@"����������̍qSU-p��iW
�2�UUR�+s�p
�H���C��B�̳,�0j
@�hIbg229ӧN�����������������������������������������������������������Ù��&hRZ���Y��8Y���,�,�P�?��霬R����T�Ђ)r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.J�U��������\i*�a\�`eUT0V���p���·-����,�0j
@�hIbg-�������������������������������������������������������������N�,�ȶX���H �,�0 ���:,$�2������*EnX*���Pga�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r��)Y ��9�V������2�T��-pʪ�cJWʐY�����:g�S��,�H�	,L�ِXXp�N���������������������������������������������������������t�p��##9bf��P �,�0 I����d��� F�2�X���j��Q9�9��r�˗.\�r�˗.\�r�˗.\�r�˗.\�sS)Y ���2�w�������q@�UUUCP��j-����t�$�e��Y�`�3BK9l��,8p�N����������������������������������������������������������:t8p�fE��$����r���,������t�VqȎD X*�P �dЂ(E.\�r�˗.\�r�˗.\�r�˗.\�r�˗8d*��IX;������l��,2���s��$��9����r�Ij,�3��,��f��&s## �Ç:w;���������������������������������������������������������Ç23�! p� Y��( �3���������Ij,B��iUUA�Uc.\�r�˗.\�r�˗.\�r�˗.\�r�˗8d*�J�������3J�p��UUR��3�rBC���:�f����9NR� Z��hIb[-������������������������������������������������������������������̋fr��� ��,�i�������w9 (eUNr�i�a�8˗.\�r�˗.\�r�˗.\�r�˗.\#C�V@"�c�������̀�$��Z�Ϊ��XC5Mq�g����s9� ,�S��,�H�	,KfFAaÇ:vvw���������������������������������������������������������·d[,BL�9j,�3��
K�������3N�ꪦ�-d��E.\�r�˗.\�r�˗.\�r�˗.\�s�V@"�c�������t�)+��*攰T��|��J�P  [���ӦFp8 �9NR̳ �9�X�̌�Ç:t�������������������������������������������������������������N�8Y�l�	� ��,�09l?������ �Wj����4EHa�r�˗.\�r�˗.\�r�˗.\�s�V@"�`$��������f
�_4��SJp�L#g��'�����Ν2	
@��Y�`���В��d9ӧN�������������������������������������������������������������N�d[,K4Z���Y��#����r�l9���8*F��UUJ��4�.\�r�˗.\�r�˗.\�r�˗8d*��IX;����Ι�S\p��UT1W9%�9frB)2���t9l$�g)�r� �f��%�l��,8s�N�����������������������������������������������������������vt�p�afE�8I���̳9K2�X�������  �����3\q�3�UT� ���ÚK�.\�r�˗.\�r�˗.\�p�Y ���2�w����f���p�!`���Ã	���΅���fr��� ��А���[2t�ӧ�����������������������������������������������������������t�p�fFE��$�2��,��p��Ζ�+`�a%�����9X8�\Ҫ��P"�0�\�r�˗.\�r�˗.\�r��Y ���2�w����l)+��J����XC�r����΅�����9K0j-FhHI��[2�ӳ�������������������������������������������������������������;:t8p�e�9bf��P �,�0 HY���Z�P�@�C��-E�����8I^
�[�
��j3�2�˗.\�r�˗.\�r�˗8d*�8������[-@AȊ��,UR�4�� ����2,B�̳9NR� Z��4$$�[-��ӧg����������������������������������������������������������������̋fp�4)-@̳,��p��:t9l$��)fY�g)�r���������pʘeUP�DӜÚK�.\�r�˗.\�r�˗8dUJ�����9l�٪�(eUS�������g����Z�2��,�0j��%���dd8s�N�;�������������������������������������������������������������ӡÅ���8R  e� g-�̌�e��Z��f  ��Z� ��,�il���t�r�@0UUB Z�Yr�˗.\�r�˗.\�F� ��EP�IX;���$�C�V�v�����R39�����s4�g)�Y�`�3BBL�# �Ý:w��������������������������������������������������������������Ç2-���8R ,�2̳ ����� ,�0  � s4��  �9NR�dw��W��W��UU3&��*C.\�r�˗.\�r�˄R�Np$�����)9' �����s�P
p������в�� g)fY�PR3BK9l��8p�g�������������������������������������������������������������Ν:t8s#"ٜ�3@�Ij e�fr���fY�Qj��%�bX�!&h)-E��r�aI�,���)��
�����9�e˗.\�r�˗.\����%`���:[-E�q@SJUU,
�p�Lw���s"� 9NR̳ �9�X��fAaaÝ:vw���������������������������������������������������������������:8XY�l�f���Ij     j
@�hIbg-��fr����fY��4����[,��iNuUP����hG �r�˗.\�p�Y �����w��� 
�_�uUT�4��+�_���s"�),�R̳,�H�	,L�# ��Ç;�����������������������������������������������������������������ӡÇ2-���4
B��f��%�l�dd,,�ȶg	3B��Y�g)fZ�B����K�qJ����@h��a�r�˗.\��+ T�J���·3���ᕸUT�+�Hp�q�X����t9l$ Y��)f  �9�X��fAaÇt�����������������������������������������������������������������N�d[3���������[228p��̌��H� 2��,��s���p8T�ܰUUfMA�8C.\�r�˗8d*�IX;���'$�enX*�����T�!fg����s9� 9NS��,�H�	,L� ��Ç:vw����������������������������������������������������������������N�8XY��l�[-��fAaÇt�ӧC�d[3�&h� 2̳,�����ȳ5�Uꪦ�Q-d�E.\"�.\���	+��RZg	*e����R�r   [;����Y�� �r�e�j
@�hI��d9ӧN�����������������������������������������������������������������s�N�,,,,,,,,,9ӧN��N�,ȶg,B@�H �9K0�dw��:[+U�*���*F�p�.\���s�%`���8 8E\Ҝꪩ`T�ÄZaI�����"� 9NS��  P$$�[29ӹ������������������������������������������������������������������Ν8p�Ç���Ν:8p�"ٜ$���fY�aIbw��ZeH���UU3&��8C�˜Y ��8V?�3�a�+p,2��b��䄅�����s ��Y��)fY�Pf�&rِXXp�N���������������������������������������������������������������������ӳ�yӿ��ӡ��̋e�I� g)f �Ý����pʘeUSX����Њ\ed*�IX;��J��8f���uUT��9BB���Ö��fr�e�  Z��4$$�[29ӿ�������������������������������������������������������������������������:t�p�ae��b
@�fY��#����9� �JUT  �����g0*�J��,W���B�UUJ�!����	����Y� ,�S�� ��f��&r�l,8p�N��������������������������������������������������������������������w����t����̋fp�4Z�)�Y���#���p��p��]���d�3��P�|-���R�*��UUM)W*A�-����ȱ�e��Y�`���&r�l��8p�N�;;����������������������������������������������������������������������s�C�2-�!&h Y��)f�Ý��Å!�4����b��B�U4��
�_�uUT�*��p���dw�����@��r��� �&hIbg-�̃��ӧ�������������������������������������������������������������������������Ù��I�Z� �� ������"�
��2�����@Wa�UR���S�rLг���Ö�KQfr���f -AI�X��fAaÇ:t�������������������������������������������������������������������������N�8XYl�		��fr�` �#���rĬ"�Wj��������8�X	2;�����4 Y��)f   s4$�3���Ç:t�������������������������������������������������������������������������:t�p�����H) g)�Y���9���8�EH�
�������[�3\r�����t,� g)�Y� �f��&r�XXp�N��������������������������������������������������������������������������:t�p�"ٜ�	3KP �9NP ����f��0ʪ����Y_*F��3����tȱ�3��  P�		3��fAaÇ:w�������������������������������������������������������������������������C�2-��B@� Y��( $����������UUUT1�*�H" ����[	
K3��,�  �f��%�l��,8p�N��������������������������������������������������������������������������N�8Y�l�f�%��,�R̵!g���%�T��UUU,
���"������rٚZ�3��,�2���%�b[-��t�����������������������������������������������������������������������������N�ddg,B@�H �9NR�gw��2-A�2�UT�*�0��I�dw���e�4 Y��)f   s4�3�̌�Çt����������������������������������������������������������������������������N�d[3�&h� 2̳,�� ������ �JT�4�
�����Ι r̳9NR� Z��4$�3��̂Ç�����������������������������������������������������������������������������:8Yl�X���Y�g)fZ�L����BNI�+攰���㔱���9�HRY�g)fY�P�		,KfAaÇ:w�����������������������������������������������������������������������������p��̋fr�$��̳9K0��w����8A�-�����Z�3��,�2���А�9l,,8p�N�;;���������������������������������������������������������������������������:t�p�fE�9b
@�fY������H$�����C��KQfr�e� � s4$�3���Çt������������������������������������������������������������������������������C�dd[3���Ij g)� 	2;������:�,�3��,��	,L�s# ��Ý:t�����������������������������������������������������������������������������:t8p��"ٜ$�
KQfY�e�j3��������$� S��,��f��&rّ�Xp�Ý;�����������������������������������������������������������������������������ӧN�,ȶX���P �,�P ������[	-E���)f 
@�hIb[-��9ӳ������������������������������������������������������������������������������Ν9�l�X��%� Y��� $�?�����a ��9K2� ��BKّ�Xp�Ν���������������������������������������������������������������������������������p��̋fp�4)-@��9KQbw���:t,� g)�Y�e�)��%�l�,8p�Ν�������������������������������������������������������������������������������;:t�p�fFFr�$�
@�fY�aI�?���B�� Y���f -AH�	3�̂Çt���������������������������������������������������������������������������������Ν:8XY���3@� Y��� �-����A r̳9K2� Z��8HIb[29ӳ��������������������������������������������������������������������������������s�Ç2-�!&h�e��r���#����fij,�3��  P�	,L�# ��Ν:t���������������������������������������������������������������������������������N�,��X���Y�g)f3����C���fr��� ���hIbg-��t���������������������������������������������������������������������������������������̋fp�4Z��fY� �p��N���dg3@)�r�`�3BBL�rِXXp�N�����������������������������������������������������������������������������������ӧC�22-���9j e�f 
L�9l�ȶ[,L�� 9NS�� �9�X��fFAaÇ:vt�����������������������������������������������������������������������������������gC�d[-��L�9j  2�   ��Z�P �,�R�  -AH$�3�̂�Ç:t������������������������������������������������������������������������������������N�d[-��L�9j-E�  ,�2̳,�    � s4$�-����������������������������������������������������������������������������������������ӡÅ��fr�$�3@�HR�!Ij
B�8�		,KfFAaaÝ�;�����������������������������������������������������������������������������������N�9��l�g,BBBBBBBBBBK��[-����ӿ�����������������������������������������������������������������������������������t�p��̌�e�ٜ�g3����l�,,8p�������������������������������������������������������������������������������������������Ç22228p�N��������������������������������������������������������������������������������������Ν8p�Ç8p�Ý:t�;�������������������������������������������������������������������������������������NΝ:t�ӧN�:t�t���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������