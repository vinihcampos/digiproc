3921
500
355
1
1 1
3 0111111
139 011111011111
140 011111011110
207 0111110111011111
232 0111110111011110
235 0111110111011101
244 0111110111011100
247 011111011101101
199 011111011101100
155 0111110111010
141 011111011100
114 0111110110
30 011111010
16 01111100
74 01111011
54 011110101
62 011110100
52 011110011
119 0111100101
216 011110010011111
219 01111001001111011
237 01111001001111010
230 0111100100111100
240 01111001001110111
250 01111001001110110
233 0111100100111010
218 0111100100111001
227 0111100100111000
196 011110010011011
200 011110010011010
236 0111100100110011
206 0111100100110010
201 011110010011000
178 01111001001011
179 01111001001010
161 0111100100100
143 011110010001
190 01111001000011
228 011110010000101
205 011110010000100
181 01111001000001
212 0111100100000011
213 0111100100000010
229 0111100100000001
249 0111100100000000
61 011110001
44 011110000
46 011101111
53 011101110
118 0111011011
132 01110110101
144 011101101001
186 011101101000111
224 0111011010001101
242 01110110100011001
215 01110110100011000
187 011101101000101
189 011101101000100
157 0111011010000
65 011101100
75 01110101
43 011101001
108 011101000
73 01110011
67 011100101
122 0111001001
148 011100100011
150 011100100010
149 011100100001
166 0111001000001
163 0111001000000
106 01110001
59 011100001
120 0111000001
121 0111000000
85 01101111
78 01101110
103 01101101
68 011011001
66 011011000
102 01101011
77 01101010
9 0110100
76 01100111
17 01100110
5 0110010
19 01100011
94 01100010
123 0110000111
125 0110000110
126 0110000101
135 01100001001
147 011000010001
241 011000010000111
203 011000010000110
210 011000010000101
211 011000010000100
208 011000010000011
238 0110000100000101
239 0110000100000100
204 011000010000001
198 0110000100000001
234 0110000100000000
80 01100000
184 01011111111111
175 01011111111110
165 0101111111110
180 01011111111011
185 01011111111010
169 0101111111100
134 01011111110
173 0101111110111
245 01011111101101
197 010111111011001
214 010111111011000
162 0101111110101
217 010111111010011
223 010111111010010
194 01011111101000
133 01011111100
110 010111110
81 01011110
82 01011101
0 01011100
7 0101101
6 0101100
18 01010111
88 01010110
87 01010101
21 01010100
22 01010011
71 01010010
104 01010001
83 01010000
8 0100111
79 01001101
101 01001100
86 01001011
111 010010101
127 0100101001
136 01001010001
146 010010100001
152 010010100000
93 01001001
20 01001000
2 0100011
84 01000101
72 01000100
10 0100001
95 01000001
90 01000000
23 00111111
97 00111110
24 00111101
96 00111100
11 0011101
27 00111001
91 00111000
128 0011011111
220 001101111011111
221 001101111011110
248 00110111101110
167 0011011110110
159 001101111010
243 001101111001111
193 001101111001110
226 001101111001101
231 001101111001100
222 001101111001011
225 001101111001010
182 00110111100100
153 001101111000
151 001101110111
170 0011011101101
171 0011011101100
142 00110111010
137 00110111001
177 0011011100011
168 0011011100010
154 001101110000
98 00110110
89 00110101
99 00110100
105 00110011
92 00110010
25 00110001
107 00110000
26 00101111
100 00101110
69 00101101
63 00101100
12 0010101
70 00101001
109 001010001
113 001010000
14 0010011
29 00100101
112 001001001
129 0010010001
138 00100100001
195 00100100000111
188 00100100000110
174 0010010000010
156 001001000000
28 00100011
31 00100010
15 0010000
4 000111
130 0001101111
145 00011011101
158 000110111001
246 0001101110001
172 0001101110000
115 000110110
64 00011010
36 00011001
49 00011000
50 00010111
55 00010110
32 00010101
51 00010100
13 0001001
37 00010001
116 000100001
131 0001000001
183 0001000000111
191 00010000001101
192 00010000001100
164 000100000010
160 000100000001
176 0001000000001
209 00010000000001
202 00010000000000
38 00001111
57 00001110
47 00001101
58 00001100
33 00001011
42 00001010
56 00001001
45 00001000
35 00000111
124 000001101
117 000001100
41 00000101
39 00000100
34 00000011
48 00000010
40 00000001
60 00000000
viniciusl���������)"""9�������������������������������������������������������"9���""""9KT�����������������������������������K\���R�R���������������������������������������Ғ�������������������������������%%%%%%%%%%%%%%$DDDDDDDDDDDDDDDDE%%%$DDDG���74DDFvvvw�5"������������������������������������������e��l�[-�Õ��l�\���e��l�[-��������������Ғ���������+���l�KKKKKKKKKKKKKKKKKKJJJJJJJJJT���������������������������������������������������������������]]]]]]]]]]]]]]]]]]]KKKKJJT��T��������������������������������������������������������������ڛ��Ԕ������������������\�Ԕ���JJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJKKKKKKKKJJJJJJJJJJJJJJJJJJJJJJJJT�����������������������������^����������\ԊKKKKKKKKJJJJJJJJKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK\���ike��---------------------)))--------l�[-������������Ғ����������������%%%%%%$DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG7777777777777777������������������������WWWWWWWWWWWWWWWWWWWR��Ғ��%%%%$DDG7777777777����������������������������������������WW��777777777776��w�E%'77777774DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDE%%%%%%%"֦��e���IIIIIIIIIIIIIIIH������������������������IIIIIIIIIIIIIIIIIIIIIIIIIIIIIIII�������������������͝�����H��������������������������������������������������ZZRRZZ�---------------------)))-------------)))--------))))))))RRRRRRRRRRRRRRRRDDDDDDDDssssssssssssssssDDDDDDDDssssssss{{{{{{{{{{{{{{{{{{{{{{{{uuuuuuuugggggggggggggggggggg--)))RRRRRDDDsssssssssss{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{uuu{{ssssss{{{{{DR)RD{{sssssssssssssssssssssssssssssssssDDDDDDDDDDDDDDDDDDDDDDDD{uRr�T�^Ԕ���������������JJJJJJJJJJJJJJJT��������������������������������������������������������������������]Y�ڙ���]]^ښ���\�
T��������JJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJKKKKKKKKKKJT��KKKKKKKKKKKKKKKKKKKKKKJJT��JJJJJJJJJJJT���
JJJJJJJJJJJJJJJT��������������������������������������������������������]]]]]]]]]]]]]]]Y����������������������������JJT��������������������������������������������������������]]^��������]Y���Ԕ��]\��������������������������������������������������T����[���������������������������������������������������������������������������������]Y�ښ����������ښ��������������JJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJT��JJJJJJJJJKKKKKKKKKKJJJT���JJJJJJJJT���
JJJJJJJT���������������������������������������������������������]]]]]]]]]]]]]]]]]]]]]]Z����������������������������JT����������������]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]Y��]]^������Yښ��T��Y�Ԟ������������������������������������������������[,����TDDDDDDDDDDDDDDDDDDDDDDDE%%%%%%%$DDDDDDDDDDDDDDDG7777777777777777������������������������WWWWWWWVvvvvvvvv������������榦����w�DDDDDDDDDE%%%%%%%"����������������������������������$DE"������������������Ғ��%%$B���������%%$DDG2��������%%%%%%%$DDDDDDDG777777777777777777777777������������������������WWWWWWWWWWWWWWWWWWWWWWWV������������������������������%$DDDDG7777���WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWVvvwWWW��7��V����$Vw6v��'WWWWWWWW������������������������777777777777777777777774B֦&&��DDDDDDDDDDDDDDDDDDDDDDDDE%%%%%%%'77777774DDDDDDDG������������������������WWWWWWWWWWWWWWWVvvvvvvvv�����������������������w�4G77777775%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%"ҕ$DE"��%%%%%%%"�����������%%$DE%%%%%%%"�%%%$DDE%%%%%%%%%%%%%%%$DDDDDDDG��������7777777777777777����������������WWWWWWWWWWWWWWWVvvvvvvvvvvvvvvvv�������榦�������������������%%$DDG77777����WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWVvvwWWW��7�Vv���Vr����w7WWWWWWWW������������������������7777777777777777777777775$G��E'4DDDDDDDDDDDDDDDG77777774DDDDDDDG77777774DDDDDDDG������������������������WWWWWWWWWWWWWWWV�������������������������������wW777777�774DDDDDDDE%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%"ҕ%%%"��%%%%%%%"�����������%%$DE%%%%%%%%%%%%%$DE%%%%%%%$DDDDDDDDDDDDDDDG��������7777777777777777����������������WWWWWWWWWWWWWWWVvvvvvvvvvvvvvvvv�������榦������������������DDDG777���7��T�vvvvvvvw6t֦��w6vvvvvvvvvvvvvvvvvvvvvvvvv����vvvvvvvvwWWWWWWWWWWWWWWWVvvvvvvvw����������������������������������������������������������������7777777777777777777777777777777777777777777��WWWWWWWWWWWWWWWWWWW�vvvvvv��������֦�������������������������6vw��vw�77777774DDDDDDDG77777774DDDDDDDG77777775%%$G7�WU%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%$DDDDDDDG77777774DDDDDDDD��DG7W77777777WWWWWWWWWWWWWWWW����WVvv��������vv���vvvvvvvvvv������������������������������������DDG777�����7�Գ�vvvvvvvw�v�vv�w�vvvvvvvv��������vvvvvvvvvt����vvvvvvvvvwWWWWWWWWWWWWWWWVvvvvvvvw��������WWWWWWWWWWWWWWWWWWWWWWWW��������������������������������777777777777777777777777777777777777777777��WWWWWWWWWWWVvvvvvvvvvvvvv������������������������������V���w�DGWW7�v��777777777777777777777774DDDDDDDG77777774DDG777��%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%$DDDDDDDG7777777777777775�4DG�W��������WWWWWWWWWWWWWWWW���WVvvv��������������vvvvvvvv���������������榦������������������77777���7WWW��t�vvvvvvvvvvwWVvvvvvvvvvvv��������vvvvvvvwVv����wVvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWW�����������������������������������������������������������WVvvvvvvvvvvvvvvvvvvvv�v�����������������TTTTTTTTU��������V���w�DGWW7����������������������������DDDDDDDG77777777���74DDDDDDDDDDE%%%%%%%$DDDDDDDDDDDDDDDDDDDDDDDG7777777777777774֧W4G7Vw��������vvvvvvvvvvvvvvvwWWWVvvv��������������֦���������������������������������������������7777����7�vwW7�����������wVvwVv榦����������������������vv���vv��������vvvvvvvvvvvvvvvv��������vvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWW����������������������������������������WWVvvv��vvvvvvvv������������������������UTTV�����������������wV���������������������������7777777777777776vwW�4DDG77777774DDDDDDDG77777777777777777777777777777777��������W�777�v�WWWWWWWVvvvvvvvvvvvvvvvwWVvv�����������������������������������������������������������777���WTG���vvv��������vvvv���������������榦������vvv��vvv��������vvvvvvvvvvvvvvvv����������������vvvvvvvvvvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWW��������WWWWWWWWWWWWWWWWVvvv���榦�����������������������TTTTV��������UUUeUUUUUUUV��������U�������d���w6vvvvvvvvvvvvvvwW������������������������vwW�4DDG77777777777777777777777777777777����������������WWWWWWWW�����Vv�vvvvvvvvvvvvvvvv��������vv�������������֦�����������������������������������������TTTW77���WWW7V������������v����v���������������榦������������������������������������������������������vvvvvvvvvvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWVvvvvvvvwWWWWWWWWWWWWWWWVvvvvvvvvvvvvvvvvvv���������������������������TTV�������UUUeUeecSSSUeeeeeeeeUUUUUUUS#TU���UTU���w6vvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWW��������WWW���77������������������������������������������������WWWWWWWW���Vvvvv�����������������������榦����������������������������������TTTW7���WWVwV���vv���������tӃ��v�������������������������榦�����������榦������������������������������vvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvv��������WWWWWWWWWWWWWWWV����������������������������������������������TV������UUUecSSSSST��eeeeeeef#��U�֥��T���V��������vvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWW����WWVwWWWWWWWW��������WWWWWWWWWWWWWWWW��������WWWWWWWVvvvvvvvwVvv��wWV�����������������������֦����������������������������������TTTTTTTTTTTW����WVvv���wW�v����������U��T��������������������������榦���������榦�����������������������������榦����������������������vvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvv��������WWWWWWWWWWWWWWWV����������������������������������������������������UUeecSST��#$eeeeeeecT�U���WT��vv���������vvvvv�vwWWWWWWWVvvvvvvvwWWWWWWWW7���Vv��WWWWWWWW��������WWWWWWWWWWWWWWWW��������WWWWWWWVvvvvvvvv�����wW��������榦�������������������������������������������������������TTTTTTTTTTTWWVvv���������������������������榦�����������������������������������������������������������������������������������榦��vvwV��������V��Vt�������������������������榦���������������������榦������������������������V���UTSSUeed��##########$���������##�SUUT���U�����������v�����榦vvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWVwVwVwVvvvvvvvvwVwVwWWWV��������vvvvvvvv���������wVv�������������TU������������TV��U�����TV���������������������Vvvv�������������������������������������������������������������������������������������������������������������������榦����vv��������V��vv������������������������榦����������������������������������������TV���UUdSSSS���##$��#######$�����������#�UeUT���TU�����������v��������vvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvwWWWWWWWWWWWWWWWWWWWWWWWV��������vvvvvvvv��������vvvvvvvv����������������������������V���������UT�cV����UUed��������������������vvv������������������������������������������������������������������������������������������������������������������������榦���������vvv������������������������榦����������������������������������������UcSS�������#$���&&&&&&&&&&&&&&&&&&$&$�#��SUeT���������������v�������榦��������������vvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvv��������vvvvvvvv������������������������������������������������������TTV���TU��������TTTTTTTT�����U��UUUeed��������������������vv�������������������������������U���������������������������������������������������������������������������榦�������������������������������������������������������������������TTT�UUcT�####$���&$���������������������&$�##�UeUT�TTTU������֦�����������������������榦��������������vvvvvvvvvvvvvvvvvvvvvvvv������������������������������������������������������������������TTV��V��STTTTTTTTTTTTTTTTVSSV�����������UUUUUUUT����������������������������������������������U����������������������������������������������������������������������������������������������������������������������������������������TTTV������ecT�##$��&$�����cccccccccccccccccccc���&###�Ued�����TTTU��������������������������������������������榦��������������������������������������������������������������������������TTTTTTTTTTTV����TV�UcT��������������������UcT�UUT�����eeeeeeeeUUUUUUUUUUUV����������������U�������������������������������������������������U���������������������������������������������������������������V�����UUUeed�$��$��$���ccccCB�����������CCCCCCCCCCcc��$��#�eUUT�����U�V����������������������������������������������������������������������������������������������������TTTTTTTV��������V��������V��������������������I�z�*�������������������������SSssrjjk����������������������������������jjjjjjjjjjj�z+j�rjjjjjjjkjjjjjjjk������������������+zZ������������K
	�񱡡�qqrbbcZbbbbbbbaqqqqqqqqqqq�����
I�������������[{z��z���������jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjksssssssrjjjjjjjk���*����ꂂ�**********ZZZZZZZ[{{zZZ���********����������������@��YAA�Y%%$��� �������������������թ���5555������������������������55��yyuuyyyyyyyyyyyyyyyyyyyyyyyy��������������������������������������������������������y���555555555555A-��5y��55555555����������������55555555����������������yyyyyyyyuuuuuuuuuuA-UYYX��� ���%�����и���11������������1111111110�������$�������YYYUY--YYU�����������������5555555555555555555555555555555555555555��������55555555yyyyyyyy��������yyyyyyyyAuA�-�uuAAA--------��--UUUUYYYUU--�UUUUUUUUUUUUUUUUyAT���� �� �YYUT�������������������չ555���y����yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyAu�5�yyyyyyyyyyAAu�55�yyyyyyyy��5�u�XՁ�����������������������������������������������uuuuuuuuyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyu�Ay�uuuAAAuA�-UX� �������%%��������й11���ED�����������EEE���������0������������� �YX���YYUUU���AAAAAAuuyyyyyyyyyyuyyy���5��������5���yyyuyyyyyyyy���������yuAAuy�yyyyyyyyyyyyyyyyyyyyyyyyuuuuuuuuAAA������-----------�---UUUYUUUUUUUUYYYYYYYYUUUUUUUT�������� ����5555��yy����yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy5yuuyyA�uuuuuuuuuuyyyyyyyyyyyyyy����u-U������������������������������������������������uuuuuuuuyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyuuuuuuuuuu�AuyuuAAAAA�UX���������%%%��������й1����ED���������������EE���EE���0��������$��� �� ���YYYU--���AAAuuuuuuuuuuuuuuyy��������������yyuuuuuuuuuuuyyyyyyyyyyyyyyyyyyyyyyyyuuuuuuuuuuuuuuuuuuuuuuuuAA��������--UU-----------UUUYYYYYYYYYYYYYYYYYYUUUUUUUT�������� �������� �����������၁����yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy5�uAA,�uuuuuuuuy5y-yyyyyyyyyuuyyyA�yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyuuuuuuuuyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyuuuuuuuuuuuuuuuuA�uuAAAA���-T�� ����%%%�������и�1����D�������t:�C���00qqq33333QQmkLL.446><<AbbI288@@@@@@55VVUKKKooooooEEEPPPEEEEEEEEPP]]]^^^^^^^^^^^^^^]]]PP]]]]]]]]]]]]]]]]P]^``^]P]]]]]]]]]]]]]]]]]]]]]]]]PPPPPPPPEEEooKKKooKKKUUUUUUUUUUUKUUUVVVVVVVVVVVV55555555VVVVVVVV@@@@@@@@888888888888888888888888888888888888`````^^^^^^^^^^^]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]^]EEEEKV]]]]]]]]o^M^U@K^^^^^^^^^oE]^^^]]^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]PPEEEEEEPEEEoooKooKU5@88IIIIbbAA<<>>64..LLkmQQ33qq0tJ+���|�_/����D�Qt:\L�T[[S����PX�L���U��UUR��������QQ[��������QQTWWWWWWWWWWWWWTQQQQQQQQQQTT��TQQQQQQQQQQQQQQQQQQQQQQQ[������UR���UU�����������UU���MMMMMMMMMMMMMMMMMMMMMMMMMMN�����������������������WW����WWW�WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWQ[�[�T�דW�PWW���������TW���W�����������������������������������������WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWTQQQQ[��QQ[�������UMP�����PPO�����TTL�\L��*�$�I$�I$�I$�I)T�U|�_]�35ֶ����CC���$����###���SSUeeUUUUUT�����UUUUUUUV���TTUTTTTTTTUTTV��������������������UV�TTTTTTTV����������������������������UUUeUUUeecSUeeeeeeeeeecST��������###############$��������#######$��������###&��������������������������������������������T��������V�����������U������������������������������������������������������������������������������������������������������TTTT�cV�����UUUUcT�$�$�����CB��ƶ��37C��Q_/����A�}��a��l6�gؠP(I$�����00qqQQmmkL..466><AAAbbIII222@@@555VVVVVUUUKKUUUUUUUUKKKKoooEooooooooEoooKKKKKKKKKKKKUUUUUUUUoKUVVUKoooooooooKKKKKKKKKKKKKKKKUUUUUUUUKKUUVVVVVVVV555@55555555555@@@88@@@@@@@@888888882222222222222222IIIIIIIIbbbbbbbbIIIIIIIIbbbbbbbb2222``^^]]]]]]PPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPP]PoEP]PoPPPPPPPPEEPPP]]]]]]]]]]]PP]^^]PE]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]PPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPoEEPEU58KKKKUUVVV5@82Ibb<<<>>>66..LkmmQQ000tW��$�I(>�a��B!�D"�B6�g��(%R��E�``fff���֘\\hl||xx����Ē��ppp��jjjjjj��������������������ޖ��������ޖ�������������������������������������������������������������������jj��jjj�����������jj��ppppppppppppdddddddd�����������������������������������������������Ē��������������������������������������������������������������������ޖ��������������������޺��������������������������������������������������������������������������������������������������������ޠ����d��������jj�pd�Ăxx||llll����ڢff`�tW�T�$�P(>�a���`0�D#a���$�R�⋡��qq3QQmkk...46>><AAAbbbII2888@@@5@@55VVVVUUUUUUUUVVUUUKKKKKKKKKKKKKKUUUVVUUUUUUUUVVVVVVVVPU2<<2UPUUUUUUUUUUUUUUUUUUUUUUUUVVVVVVVVUUVVV555V555@@@8@@@@@@@@@@@888228888888822222222IIIIIIIIIIIIIIIIbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbIIII]]]]]]PPPPPPEEEEPPPPPPPPPPPPPPPPEEEEEEEEEEEEEEEE@qA^KIo^EEEEEEEEEEPEPEPEPEPEPEPPooEEPPPP]]]]]]]]PPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPEoU5@EEEEEEEEEoEoEoEoEoEoEoEoooEoooooEEEEooKKooKKKUUUVV555@@@222IbAA<AA<>6..LkkmQq0t:��T�P}�a��B���8.��.��n۶��ϰ�B6}�)U��|�(�L�T[Z�������X��RRRL���MU��ՐQU������������������������UUU���MMMMMMMMMMMMMMMMMMMMMMMMMU�������������������MPRRRRRRRL��������RRRRRRRL�RRX�����RRRRPPPX��RRX��������RRRWWWWWWTQQQTQQQQQQQQQQQQQQQM�̑M[�W�QQQQQQQT��QTWWWWWWWTQT[�U�QQQQQQQ[������������������������QQ[���������UUU�MMP��X�PO����[[[TL�L�E|�(>�a�����,;ð�;ð���8/+����ؠIJ�R�⋠���E���10�����������%%$�������� ����������������YYYYYYYYYYYYYYYYUUYYX�������������������������������������������YX�� ����������������%%%%%%%%%%%%%%%%%%%%%%%%%%%�����������������������%%���%%������������uuuuuuAAAAAA�A5A�@�AAAAAAAAAAAAAAAA��AAAAuuuuuuuuAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA�-X�����������������--����������---U-UUUYYX� ����%%����й1��D��ED���Q_/��RIA��A����K�)JR��)JR���04ù.��`���(	)T�E�`�⢢�֘�\\hhl|xx����Ē�ddddddppp��pdd���p�jjjjjjjjjjjjjjjjjjjjjjjj����jj��������������������������jjjjjjjjjjjjjjjjjjj��ppppppppppppppppppppppppppp�����������������������Ē��Ă���xxxxxxxxxxxxxxxxhlx�����xxx����Ă����������Ġ�����������������������������������������������p�����ܚ�������������������������ފ��������������������������������������������������������������ފ�ޖ�������������������������ޖ��������ޖ���������jj��pppddd���Ăx||ll\\���ff�f�`�(�����A�����p%�a�T�)$ID�$ID�7Ҕ��a����p�!�JU|Qt������& ��11$������ *�� �       �������������������                     $��������11111111111111111 ��� � �� ��� ����((((((("������������������������������������������/.�.�((((((("��������������������((((((((((("���������������������������������������������������������������������������������������������++���  $��11 �&6����:
)RI@�!����p�h5�aM�Do�ADAID�JXV�a��;��8/+��b�U|Q(���������& ��11111$��� ��$�                ��   $�$����������������1111111 ��������1111111 ��� �� �"�������������������������������������������������%�%�%Ȩ��������������訨�������訪


��������������������������������������������������������m����im��������iiiiiiiiiiiiiiiiiiiiiiij����Ʀ��FFI),LLH(('���ƅ�Ɇ�ɍm�&n.���*I(>�gm�y\%��R���$F�گ�����_��~/�A��D�JR��a�w%�p\`�l�	)U񁁃����k[[Zaq�������

JJJI���	���������������������������������������������������������������������������JJJJJJJJJJJK














	���������������������������񱱱������������������*******+{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{zZ�+�ZZZZZZZZ[{{{{{{{{{{{{{{{{{z**����*******+{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{z��{{{{zZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�������������JK
	���񱱡rbbc[[j�����|�J�Ja���p\%���)"H���_�����rnMɹ7&�ܰ����v��o�,+aܗ�Fϱ@�It:L��[[Z�������PPPPPX���RO�[PŘ�������������������������RRRRRRRRRRRRRRRRRRRRRRRRRL�������������������RRX��������������������������PPPPPPPOPPPPPPPO��������������������������������������������QQQQQQQ[����������������������������������������W��TQR��������������������������QTQQQQQQQ[�����������������������������������������������ՕR��������������UUUUUUUUUUUUUUUUUUUUUUUU���MMP��RRRX�PPO������TL�]��|�$�a���8Ka�T�o�j�K	J/��ϼ�ϼ�ϼ�Ą�����XJ�_ĉ����05�r]�l!>�ID��0qq33QQmkLL..>>>><<AA<AAAbbbI.b2._/���RRRRRRRL������������������RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRL��RRX���������������������������PPPPPPPOPPPPPPPO�������������������������������������������QQQQQ[������QQQ[��������R�N�[�������������������������UU�MU�U[��������QQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQ[���������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUMMMMP���RRRRRX��PPO���������[T\]��T�I(�����.�%#x��W��a)D����>��>��>��>��>��>�������_��A����a��y]��l�J��&&fffj-�e�ƅ�Ɔ������Ǉ��(((((,LI)))))))))),LLLLLLLGI,G���))))))),LLLLLLLH((((((('�((,LLI,LLLLLLLI)))))))'	'ƅ��),LLLLLLLH((((((('��������������������������������������Ɔ�����������������������Ɔ��������������������������������������������������������iiiiiiiiiiiiiiiij����ʩm����������������������������������������������������������������iiiiiiij��������j������������������������������Ʀ��FFI)),I),LH((('����Ɔ����ɍm��*..�A��E*I(>�c���aM�گĢnI��7O"7F���tn�Ѻ�.��/���ܥ�����H�,+
�.��#bJU|Qt8������� ������1$����������1111111$��$��������1111111 �������� ��11111111111111111111 �11111111 ��������7�����������������������������%��������������������������������������������������������������������������������������������������������������������������������������������������   $��11111 ��&&5������J.�B��P}���m�p���{�_�%��}��Ӵ�ԡa"r'"r'"r'"r'!r6��n�q���Qa+�A$M��ù.��$�JU|Qt8������ ��111111111111111111$� �11111111 �������� ���11 ��������1111111$� ���������7������������������������������������������������������������������������������������������������������������������������������������������������+++++++++++++++                  $���11 �����&5�����������E*PA�ۂ�0�;�{�a)Dܾ���iJr!7�x7�x7�x7�xJwr'#a��/"�ϼHR��F�E�aA�;��`�ؠIJ��.�ִ������CCCCCccc���������&&&&&&&$��&$��&&&&&&&#�������������������&#��������$�ccc����������������������������������cccccccccccccccc�cccCCCCCCCCCCCCCCCCCCCCCCCCCCCB��������CCCCCCCCCCCD����������������������������������������UUUUUUUUUUUUUUUTV��UT��T����������������������������������������������������������������UUUUUUUUeeeeeeeeeeeeeeecSSSSSSSS������������������##$���&&&$��������cCB��������7B��IJ�J``1�p\��%&���XI�}��}�t�#u�܈�Ҁ�	 �	 �	 �	 ��(��XE(R��^E�}(��j �&�
r\m�>ϱ%*�(�]&j-�mi�����Ɔ������������Ǉ��((((((((((((((((,H(((('��((((((('�������Ǉ��������Ǉ��(('�������Ǉ�������'���������������������������������������������������������Ɔ���Ɔ������������������������������Ɔ�����������iiiiiiiiiiiiiiiiiiiiiiiiiiiij��ʪ������������������������j����mꪪ������iiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiij�������������������������������Ʀ�������FFFFFFFFFFFFFFFFFFI),LLLH(('��������������ɉ�mmj*&n.&�AE*P(I/���y\�a�Vo]�	7/�����]�(\�����D�oF�oF�oF�oF��@}Ѹ%�9���I�}������7��+�<�؄B6}�)U����0q3QmkkLLL...4...444666666>><<<<<<<<<<AAAAAAAA<<<<AAAA<<<<<<<<>>>>>>>>>>>>>>>>>>><<<AA>>>>>>>>>>>>>>>>>>>>>664>>>>>>>>66666666>>>>>>>>66666666444444444444444466444...............................................KKKKKKKKKKKKKKKKKKKKKKKKUUKKKU55UUUUUUUUVVVVVVVVVVVVVVVVKUVVVVUKUUUUUUUUKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKUUUUUUUUUUUUUUUUVVVVVVVVVVVVVVVV@@@@@@@@22222222IIIIIIIIIIIIIIII2IIIbbbAAAA<<>>>>>>66644LLLLkkmm33qq0tJ+�K��
`c��85�JM�گ����.��nBn��H��E������<���7$���p7�"rv��$,%/�j7�,3�༠���(R�R�E�`f����֘��\\\��\\\hhhhhlll|||||||||||xxxxxxxx|xxxx���||||||||llllllll||||||||||||xx��llllllll||||||||l||x|lh\llllllllhhhhhhhhllllllllllllllllhhhhhhhhhhhhhhhhlhhh\\\�\\\\\\\\\\\\\\\\\\\\\\\\��������\\\\\\\\\\\\������������������������������j����������������������������jj������������������������������������������������������������������������������������������������������������������Ē����Ă���xx||||||lllhhh��������f��`�(�J+�K��
`c��9,;���_�$ܾ�v��n�@��h���{����7����oe��H #r�@Jwr1�n�}(����}�r\���bI%*Q(�L�[Z������������������������PPO����������������������������M�����������������������������������������������������������������������������������������������������UUR����UUUUUUUU��������������������������������UUUUUUUR������������������������UUUUUUUU��������U�������MMMMMMMMMMMP���RRPPPPPPPPPPPPPPPPPPPPPPPPX��PPO����������TL��\L����J�a1�8,85�aIj�M�ia!r#w7�7�_��W�n�v�np_���oc{��+�r�����NF�.�����Ҋ�F�}�r^Wl!}�	T�%*�(�L�T[[[Z�������������������������������������������������������������������������������������������������������������������������UUR���UUUUUUUU��������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����������������MMMMMMMMMMP���RRX�PPPPPPPOPPPPPPPPPPPO����������TTL��\L��|�J�_a�1�yA��0�H޿�!}�t7\�Ȓ��Cr�G �Mڿu����M�n3q��np7a�M��_�ܾ�(����$/�nW�� �,3�༮؄lP$�I)T�E�`�⢢�����֘�������hhhhhhhhllllllllllllllllllllllllhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhh\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\������������������������\\\\\\\\��������\\\\�j�j��������������������������������������������������������������������������������������������������������������������������������pppdddddddddddd�����xxxxxxxxxxxxxxxxxxxxxxxx��xxx|||llllhh\\\\\\�������ڢff�``�tW��$����ۂ༮ 5�JM��}�ia"7�p7����F���^Jy�y���� w���n5���n�{9�rn	@�L"�/����;Q�aXw�yA�gؠI$�R�⋠����EE�������������������������������������������������������������������������������������������и���������������11111110��������������������������������1111111111111111111111111111111111111111111111111110������YYYYYYYYYX���YYYUUYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYUUUUUUUUUUUUUUUUUUUUUUUUYYYYYYYYYYYYYYYX��������YYYYYYYY ������%%%%%%%%%%%��������������������������������������и��0��11�������D�������(���RIA���r\�7��~%�}�J"7�@v���nѸ@+����ӴRA�Cy�2A�_�@��/�n2A���_�ܾ���(MѺ}������\��v��gؠP(R�A���������kkkkkkkkjbbbbbbba������������������������qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqrbbbbbbbbbbbbbbbbbbbbbbbaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqrbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbc[[[[[[[Zbbbb��������������������������������������������������������������������������������������������������������������������JJJJJJJJJJK
	���������񱱱���������������񱱱����qqrbbbbc[[[kkkj���������Q_%R��K�6�W�r\�i�H��
�7/�n�됥 Ѐ�����k���H3�b�e~�ɵ�y�#�U��A7��ؿ� ��nI ��n���������0�K��b���>�J���t8������������������������&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&5����������������&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&5��������&&&      ����������   ���������������������������������������������������+++++++++++++++++++++++����������������       $��11111111111 ���&&5����������������:��*�$�
��B��ð�)" �+�(���v�7w���\������y�v�o9~��� B<�a�a�b���k�<������_��W��Sz}ѻ�����!J,%~�H5�r\�!��b�%*�(�L\L���TTTTTTTZ������������������������������������������������������������������������������������������������������������MMMMMMMMMPMMMMMMMU������������������������MMMMMMMP���������RRX���PPPPPPPPPPPO����������[Z�[[TTTL����L���|�J�J��A�+�� Ԥov����y��i@���W�n7�W�v� i �@�ﰅy_������#��M� w�D�sq��oB7M�����}�����#a��P$���C��������������͵�������������������������������������������������������������������������������������������������������11111111111111111111111111111111��������111111111111111111111111������������������������� ����� �������� ��������YYYYYYYYYYYYYYYYYYYYYYYX�������� ��������%%%%%%%%%%%������������������������������������и��1111��������EED��������Q(���RI$��>ϳ�6<��������	$/��)B�&�7+�_�ƿ��N�$�ca ^@�O�����_���(�/&B /�0�e��K$���Q�7"J�}�r�W��o��3�/+���b�%*�(��33333336�������ֶ��������������������������������������������������������������������������������������ֶ����������������������������������������������������������������������ƶ��������������ֶ���S��$T#���#$���#���SSSSSSSST��SSSS��$��#��#���SSUeeeeecSSTd�3$��#SSSSSSSST���#%c�&$�$�$���&$������������cccb���������������������������������ƶ�����37C��Q(�W��$�P}�``1�y\%�a��H��I�}�i�Bn� �݂_��^M�  
���'+��N@^N�/�_��}~�V�&ݢ/� w���n%�/�n_toB�/�nXK�$R��aܗ�v���P$�R��C������������ED�������͵�����������������������������������������������EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE��������������������������������11111111111111111111111111111111111111111111111111111111�������������$� ��0����%%%$����� ���������� ����%%%$�� ��� �� ��YYYYYX��X���-$��������� ������Ɉ�$���%%������������������111111111111111111111110��������1������EEED���������(�J%�U*I(>ϰ��n���;o�+�����v��r'���������o! ��@^B<���_�o4�c���������a��h�{��w�M/������	�Ar��9���!a.ԑJXV�/+�F�JU*Qt:&.&fffffffffffj*******-����������������������������������������*******************************-������������������������mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmf�,LH,I,LLLLLLLI)&FFGI,LI&G����������Ʀ��
����F�FFI)'��ǆHLLH('���������������������Ɔ���ɉ�������mmmmmmmmmmmmmmmi��������mmm��**&fffn..&�C��Q(���T�$�P}��`c��.�ÃXc}گ�HM��r4�v��� ��p�+��d@����>�C��7�M簇a}�y7�������h��Ŀ�;@���_p���7�)Kr\�#gؠIJ�J%C��������������������EEEEEEEEEEEEEEEE��������EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE������������������������������������������������������������������������������������������������0��T������%$�����������������������������%��$���������� ���YX�� �������� ��Y�U ��������������%%%���$Ɉ������������������������и��11�����������������������������������EED������������tJ+����I(a��B�o+����k
H���_|�%���ܯ��&�_���ݢ�a��a�5��2��������v7��k��y�&o'',!X@��y���n�{/�ލ�Ȇ��>��_�	������p^Wl!>�I%|�(�J.�C���t8������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������&6��� ����11$������������������$��$�111$�   ����   ����  �$�� $���111$� ��6��&&&5���������������������������������������������:�AD�Q_/��R�@���"c��.�ÃA�H޿���}�J"7z#{��o �E1�c�G�#{�'������}�os��ϻ_v�����o0���ɐ��y@#p7��F�&���
�M���a�w�p]�l!}��JU*�_J%�D��t:\\\\\\\\\\\\\\\TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTL��������������������������������TTTTTTTTTTTTTTTTTTTTTTT[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[Z������������.��CF����Cc�������&&&&&&&&&&&&&&&&#��#$�$$�$$�###########��#���ST���#����#���#######$��&&$�$f�����cccb�����������������ƶ�����33333335337C��Q(�J%��|�J�g�l!���p\%��������!}�ia"7_���P�ݢ/��`@���@C��>�/�7���n+���7h���ד�� /��@��_���� $��"�/�HXK�7����aܗ�y]�`�l�	)T�U*�_/�+�D��t:fffffffj*******&fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffj***********************-��������������������������������������������������������mmmmmmmmmmmlM��Y�kkZaq����������








���K	��JK
JI��������JI����������������J�I�JJJJJJJJK

	�����
	�[���񱱱��bbbbbbbbbbbbbbbc[[kkj�����������������������������������������������(�J+�E|�_%R�W��D �m�y^W�a��3o�,$ܾ���#r#p�/�O%/�� �!�B<��B�����n#q��F�7���n/��'sy���aH;�b7����zv�P0�Ⱦ�ﰕ�H��Kr\�vݱ��(	$�JU*�_/����D�Qt:����������������������������������������\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\L������������������������TTTTTTT[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[Z�����������Ş˟bK���kkZaq��������������������K���K


I��������JI��������������
�I�KJJJJJJJK

	���qq���r��񱱱���bbbbbbbbbbbbbbbckkkj�����������������������������������������������(�J+��D��_/��T��6A�۶������7ݫ	$/���u�܄���$�k���m�3�����A���oq���>�7���{����M���a��w��n5������xr7i7O��W�"o�,05�p��v��gؠP$�I$��U|�J����D��00000000t:�C���3333333333333333333333333333333333333333qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq333333333333333333333333QQQQQQQQmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmkkkkkkkkkkkkz��Fϱ�i��ͬ�٬��٭������������������������������%%%%%%%%�����������%%$�����������%%%���������������������1��11111110�111��������EEEEED������������������������������������������������t:�C��Q_/��T�U�}��a0�.��Xf�J]�!�F�iB�)@H F�_��k���H8� ����a���yﻏ�����7���}�7����B��y6 j��%���N@7�@7"Jt��܍�y�\��y^Wm�F�b�@�I$�R�T�U|�_J%C���t:���F�ֳCC7C���kj���Yq�kkkkkkkkkkkkkkkkkj����k[jbci��a�kkkh�X�{���*�;iV�CC5󉚉q��a���������������������������

JJJJJJJKJI��JJJJJJJJJJK




	���������񱱱���cZbbbbbbbbbbc[[[kkkkj������������������������������������������������t:�AD�Q(�J%��|�_%R��K����c��.��Xf�JF����7]��M�������by~�� �O��<��w�_�~��W�_�~��M�7�n,!�N��0�a�l@���K_��� /�7�"����ɹ��}��.���0!�I$��J�R�U��|Q(�]�C���t:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\L\\\\\\\\\\\\\\\\\\\\\\\TTTTTTTTTTTTTTTTTTTTTTTTZ��K������[M��TL�\[[[[[[[[[[[[[[[[Z��L���[J.�6�CF�����QR!QKԱ1Ġ6(:Zϋ��[S���������������������PPX�����������������PX��RRRRRRRRRRRRRX��PPPPPO����������������������������[[[[[TTL������\\L�C���t:
%�D�Q(�W��U*I$�_g�l!�m�p\$�0�)�7�V����F��ܯ��&�7��!���i���yO&f��v��}�7��ڿj�� �ń;���!M����d�_�����F��r�F�D�aA�K�༮۶�F�b�@�I$�R�T�U|�_J%C���t:���F���54�f��k[Z���kkkkkkkkkkkkkkkircj��������Y���E������x��_bJ���Ѭ���l\hhhlll|\\hhllllllllllll||xxx����������Ă�����������Ē�����������Ă��xxxxxx||lll||lllhhh�\hhh\��������������ڢ����fff������``�t:�C���t:�C���t:�C���t:�C���t:
%�D�Q(�W����|�_/��T�$�P(a��Bvݷ��p\$�0�(� �+�(���aw7�_��M��X��$��7���^L�缀�os�Ѹ��~��^@�_���o0��G�'�b���Y �� Bn	@�n��ą(����JXV�p^Wm�v�����(	$�JU*�J�W���D�Qt:�C���0000000000000000qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq000000000000000000000000qqqqqqqqqqqqqqqqqqqqqqqqQQQQQQQQQQQQQQQQQQQQQQQQ.qt(�&5�&6��(���(ؒ`�\h������������������\�֢f��fl\�fff������"J�l�%A�����l��}�������������������PPPPPPPPPPPPPPPPPOPPX���PPPPPPPPPPPO���������������[Z��[T[[[[[[[[[[[TTL������\\L�AD��t:�C��Q(�J%�D�Q(�J%�D�Q(�J%�D��_/�����|�J�R�T�U*I$�J�����`1�y^W�p�k°��ڻU��_q(\�(t "oe�������&� ������hɽ��>�}�7���n&�>�7��zy
�r��	 �!��k�7���݄^E���	_ĉ����;�༮۶��ϳ�P(I$��U*�J����D�Q(�J%�D��t:�C��````````��������������������������������````````````````````````�����������������������⢢����������������������\��QmQm.Lmq0QQ}�Q�$����1������������������1�D���̢f֢�(��(��������������X��05*�fImmmmkkLLkkkLL...4444444466>>><<<<<<<<<<<AAAAAAAA<<AAAbbbAAAAAAAA<<<<>>666666444.444...LLt��������������������������:�C��Q(�W��D�Q(�J+���|�_/�����|�_/�����|�_/�����|�_/�ĒI$�I$�I%�@��>ϰ�l!����y\�rA�3
»Wj�W�7IB�&�n��{���H;ɇ�����N�A�_�~Ѹ���k��ݣq}�a}�v�_��� ���	���A�J"a�}�����"o�,3�<�۶Fϳ�P(	$�JU*�J�W���D�Q(�J%�D�Qt:�C���00000000qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq000000000000000000000000qqqqqqqqqqqqqqqqqqqqqqqqQQQQQQQQQQQQQQQQQQQQQQQQLQ3Q0_����5���[Z��\L[[[[[[[[[[[[[[[[[TL��[Z�&��f***** � ��A�G.���<DD<\���[\L���TT[[[Z������������������������PPX���������������j-��*&fffffffj*&fn.....&�C���(�J+���|�_/�����*�J�R�T�U|�_/�����|�_/�����*�J�R�T�T�I$�I$�I$�P}�g�l6D"c����H5�aXRD�W�}��Fn� "�����v� j��� ����a a�7���7ݦ�<��a�f���F/&��;E_�F�_���P9P��B�W��$M��/+�D#gؠP(	$�JU*�J�W���D�Q_/�����|�t:�C���t:�C���qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq000000000000000000000000qqqqqqqqqqqqqqqqqqqqqqqqQQQQQQQQQQQQQQQQQQQQQQQQmkLQ$�iR�6���Cd�����7����������������75���6�G7A����茔<Td(d�x�S336���ֶ�����������ccc������������������������&#������������cccCcCCB���������ƶ�ֶ���33333333337C��QtJ%��|�_/�����|�$�I$�I$�IJ�R�T�U*�J�R�T�U*�J�R�T�U*�(
�@�P(>ϳ�6�"0���.�a�V�JIj�_}���rxv����sq����s�Ǔ%�ѯ'� �'v����7���������j�1 D a1�*�k�_������R����o���%�y]�`0B!>��@�I$�R�T�U*�_/�%��|�_/������t:�C���t:�C���������������������������������������������������������������������������������������������������������a�h��}���*&m��**-eƍ����������������*)���n�"J����ffffFFFFJ�}������������>�{634Lt>�m���-�����ɉ�mme��Ɔ���Ɔ������Ǉ����������������������Ǉ������Ɔ���ɉ��ɉ��mmm����*&fffn..&�C���(�J+���*�J�R��I$�P(
�@�P(
�@�P}�g��}�g��$�I$�I$�I}�g��}�g��}�a��l!�F�a��l6���`1�vݷ��p%��A��" �ĢH_y���M���@��H#y���}���+��{�!^O@A^N�!�C��y:y
o-��G����_��������P�����J+�AҔ���.���g��}��@�I$�R�T�U*�J�R�U��|�_/���AD��0q300000000qqqqqqqqt:�C���qqqqqqqq00000000t:�C���00000000t:�C���00000000qqqqqqqq33333333QQQQQQQQ33QQmmmmQQQQQQQQ343QA.qAQQ5mm@qqmmmmmmmm6.kmkkQ0t���������J	�I�E�D̢�|^^rFJJ�}����������@A.��Ԕ���:����S����[[[K����������������������������������������������[[[TTL����\\L�C��Q(�J+��U*�J�R��I$�P(
�@�P(
�@�P(>ϳ��>ϳ��
�@�P(>ϳ��>ϳ����a��BD"�B!���m�v�W��p%��A��" ��H_}��둥����_��Bv�H;ɧ��!O��7���y��u�u��+�j�7�7����� w�����<���ȘE�_}��Q��JXV�+�6�g��(
I$��J�R�T�U*�J�W����|�_/�����0q00000000qqqqqqqqt:�C���qqqqqqqq00000000t:�C���00000000t:�C���00000000qqqqqqqq33333333QQQQQQQQ33QQmmmmmmmmmmmm.>3t&8���΃F������������3B������asZ�����p[^T����`ھ1//9##%}>�O��興���d<DdD��D@Q$�nT��ڢ�QJ���������&&&&&5�5����������������:�C���(�J+���|�J�I$�I$�P(g��}�g��}�g��}�g��}�g����a��l6}�g��}�g����a��l6�"0�D"�B!�۶�+��8K�R�|ov�$ܾ���#7spv���n���J_��5�v<�a
�a�����F���7�oy��G��&M����q����oF��NF�&萯�o$XV�a��v��a���>��@�I$�R�T�U*�J�R�T��|�_/����E|�_/�.�33333336��������35���ֶ�������C�B���q�ED�D�x��������\�f�ff�_:
%6����A���R�h`�IQ4t%����������������������C���C���.0lIt��TTT[[[[[Z�����������������������������������������������[[TTTL���\\L�AD�Q(�J+���*�J�I$��@�P(g�����B!�D"�B!�D"�B!�D#a��l6���B!�D"�vݷl��`0�n���+��8K�R���v��(��y�r$�}ѽ��� �]����Cɦ/�� ���F��_��}~�V/&�M���Cq���B�Gh%�����Q_�y"o��05�pWl6�g��(
I$��J�R�T�U*�J�W����|�_/���U*�t:\\\\\\\L\\\\\\\L\\\\\\\\\\\\\\\L��������[[[[[[[L��T[[[[SK��Z�����K��[S�J%A��������(&53�8��O)A|A
??==1/99#99##%%%"}�������ŋ ��J��������������&&&&&&&5����������������:�AD��_/���U*I$�J�A�}��g�l6D"`0��`0��`0��`0��`0��`0vݷm�y]�m�vݷm�vݷm�y^W��p\�rXph4¥&�����$&�n��% <���$�Bv�� �M ���" ���}���A�$@�%/�ݫ�y ܾ�Ȓ��_p����7Җù.���g��}��@�I$�R�T�U*�J�R�U��|�_/�����*�J���33333336��������35�������������DƳcG2��5�f��������ƶ��C�cF��CD�2�$�P}����y�+{zTBf�FͯC�53���󓓓�222QR'��Ɉ�8��8��H�l�<�bK��`�ff�������֘���\\\hhhllllllllllllllllhhhhhhhhh\\\�����������ڢ��fff����``�t:�E|�_%R�T�$�I(
�����a�B!�A��m�vݷm�vݷm�vݷm�vݷm�y^W��y^W��vݷm�vݷm�y^W��y^W��vݷm�y^W��y^W��y^W��vݷ��y\�p\�a���k�{�a)Dܾ㴰������M�n� ���
�N��/��m�cɁ  y0�i�����;E;�K���+��@J#v��}����})JA�;��<�؄B6�g��(
I$��J�R�T�U*�J�W����|�_/�+���|Qt8������������������������8��������8���������������������������������������������������������6����S���bbbbbbba�Y����P�R�B�*I42_�ä�eY�JD%mH,QQML�������ļ��������""}>�B� ��W�Y�DP(R�⋡Т������֘��\\\hhllllllllllllllllhhhhhhhh\\\����֘������ڢ�ff����```�t:
%�E|�J�R�RI$�P(>ϳ�6��0!�۶�+��+��+��+��+��+����.��/+��+��۶�+��/+��+���������9,84��I"�W�Q7/��)B�.B��7��	 ����g��_��rA��7�o9�7h�y�A���oD�n�/"��儈$�R°���p^P`�l6�g��(
I$��J�R�T�U*�J�W����|�_/�����0q00000000qqqqqqqqqqqqqqqqqqqqqqqq00000000qqqqqqqq00000000qqqqqqqq33333333qqqqqqqq33333333qqqqqqqq33QQmmmmmmmmmmmmmm.q_1.�&_f�T��[[[[[[[[[kY��Ë����d�E����ښD�ā��@o> ���OOO���OOLLIINLLNEDNIH�EB�A@A�E����`�l�	)U��ֶ�������CCccccccccccccccccCCCCCCCB���ƶ����ƶ�����337C��Q(�W���U*�$�J�A�}��a��B!���`0�o+��+��+��+��+��.��.��.��.��.��.��o+��.��<�+��+��+��.��8.����h4�%$��_�Dܾ��"�f�H� "n#v��璍�_��A�C5�7h�����/%���F�7��W�7/�7�"�营� ��K
°�;��`��l6>ϳ�P(
�I%*�J�R�T�U*�J������|�_:
%A�������������������������������������������������������������������������������������������������������kkkj����������Y��x��6J�=L�-������������P2&�Q������do�{�!
���&��F����EEEEEEEE55555553������7�X8�xxx (s����k�J��Z�L�K��͐PM��O��͍��ˋ�����������[[[TTL���TL�L�C���J�I$�I@�P}�g��}��a�B!�۶�+��+����.��.��.K��.K��9,;�<���8+�.��8��8��8��8��8��8��.��.��8K�� ��7�j��JQ$/�n�둹��@ޗ����~��7�k���o!���<��
�o%~��r�˴��܌n���r������\��y]�`�l6>ϱ@�P(
�$��J�R�T��|�(����D��tJ%����000000000qqqqqqqq33333333qqqqqqqqqqqqqqqq33333333qqqqqqqqqqqqqqqq333qq000Q333qqq0t8��	.)�'���GA�T��I6k3kJ��
.H�Y$lPt�I%���d�x�hP���&��T�ov�����3g`3<3
|B����@�/���vbT����������������OOOOOOOLK�H�DB�`��##""!��N�Q�RĴ�5�%|�qq4<<4L.Q(�L�N������������������[[[TTL�������L����Q_%R��I@�P}�g�l6�"0vݷm�y^W��y\�p�p�p�a�v�a�v�rXv�a��K�o�ے�0���.K��.K��.K��.K��8��8��.��.����.Ka�S|ov��%r����XE�\��toK�_��n���	�q���f�7�W�$�������toD�.�n�p���7�,04�8��D#a���}��@�P(	$��T��J�W���E|�_J%C��Q(��33333333333333373333333733333333333337337G���٬�h6(���s��*ڢ�\Kz�.�<��W٩Q��m>	/6}�[��(��%*jJ�~"޼D��r�<�V�4*zbU�R�3�>*����������������zzzzzzzzzzb^rFJ�"%l����J&i���A�t6�&5��&&&&&&&&&5������������������:
%�E|�J�I%���>�a��B!��m�v�W��y\�p�p�%�a�v�a�v�a�ph4�A���JM�})a�f�rXV�pv�a�v�a�w%�r\�%�r\�%�r\�%�r\��p�p�p�%�a�pk䈂�W�	J$���Dn����P>�n^H�_�M��v��݆�7a�W�n' � @]���p7�wr1�n�y�Ҋ�v��
���༠��l6>ϱ@�P(
�$��J�R�T��|�(����D��tJ%C��������������������������������������������EEEEEEED��������������������EE��D��������͵��|Qmq5�>�E% �W`��(������H	���B���Z���$�%�:�zTB�X�2^
� T�ֈN�*�%;B�N��&TꚚ������������������������鉉yy�))+�T,T,D(4X��y�QLLe�F��d���������������ƶ����337AE|�J�R��IA��"�;n�������9.Kð�;ÃA����A��h4a�f�a�f�aR���7��})�R���M��a�f�a�`h4�A���a�v�a�w�p�p�r\�%�a�pk¥&�� �+����}Ǒv���nB���y#���r�\�� ����Sz$xJ"r#����	�_��oJX`kø��#g�l6}�b�@�P(
I%*�$�R�U��|Q_/���E��(��33333335��������35�ֶ�337A����!}�
 ǷRJ�أ`\!���mRt*���NF�%!Zchs���J����q���Y:$��Dɍ	RbD�&t�Ҥ:L�T-����������������OOOOOOOO��OLLLK�LK��NNH�IH��H�D�$dDO�RW�����xP$�M�L[[Z�����������[[TTL����\\L�AD��J�I$��A�D �`1�vݷ��y\�p�%�a�v��Xf�a�f�aXT�)JR��)JR��)JR��)JR��)aXV)JM�D�aXc|A$A��E�aXV�aXV�a�f�a�f�A��h5�r\�%�r\�%�r\�%�a�ph5�a�S|�$F����I�}��7F�(\�ȍ��N����zy"�\�� /��$y!�;@��ȘE(]��>�!J,%ڈ&�
a�v�p^Wl6>�a���
�@�P(I)T�%*�J�����|�(�J.�C���000qqqqqqqqqq33333333QQQQQQQQmmmmmmmmkkkkkkkkmmmmmmmmkkkkkkkkmmmmmmmm33QQQmmmQ333qqq0.QL�Q�� a�Lx���;	)E�Yؠ�� ]�\�%_��5�Y�bωَ�f&�����o���ɭ*�L�16��D�u�ӨZ'????????????????============111/=111////"""""""%%""}>�H�MW�Bb�%���E���1��������EED�����������t:
%�U*I(g�l!��m�y^W�p\�a�v�Xf�aXT�)JR��)7��|�$M�|�7��|�7��|�7��|�7���)JM�DAv��)a�����&��o����o��+
°�+
°�3�0�3�0�;ð�;ð�K���84��3
��&���]��a)D����;H�r7"Jx7p}� ;@ލ�ލ�ކ�n]�H��B�o"�/���儯��7�)Kù.K�༯(0B6}�a���}��@�P(	$��T��J�W���E|�_J%C���000qqqqqqqqqqqQQQQQQQQQQQQQQQQkkkkkkkkLLLLLLLLkkkkkkkkLLLLLLLLkkkkkkkkmmQQ333qQ333qqq0Q^P6m$�I)�`F����XE�_���r�U��Z�NFu�9�G� lϊ��D�*~u��ӢX�ɉT���ևN�htIӧN�BѢt-�????????????????========111111//=111///9==?SSS1/9##/?=/%//19""w��8���&j-��*********&fn...&�C��Q_/��RIA�}��a1�v�W��p\�p�$��3°�*R��&��o����H�$��7��x�7��x�7��x�7��x�7���H�#{�a)Dn��|��|o$ID�$ID�JR��)JR��)aXV�aXV��A��h4r\��a���h5�a�f�JR�Av����rH_x�;JP���������>��O�}Ѹ��%��P���}��7,%;WjH�,(5�r\�%�y]�`�l��g��(
�@�P$�R�RJU*�_/����|Q(�]�A�����������������������kkkkkkkk[[[[[[[Yqqqqqqqrbbbbbbbaqqqqqqqs[[[[[[[Zc[i����QQ333qqq02y�""�>��qxq%ԕL���^A���t*�g��&MQ�񡉊�H>��h����Y��hM�!��I6f��*�:թΓhu
t�ӭB�:s��������������������������������������茕�rJ�}���EH����_DC$O��sEE�E�`�f�ڢ�������fff���````�t:
%��*�$�g���A��m�p\�p%�rXv�a�f�JR��)7��|�$ID�$F�ADADAD�o��o����Dڰ�B��r7W��J)E���o��o���)JR��)JR��)JR��)JR�h4�A��%�a�ph4�Xf�aXVo]��_�%(�rH_q�]�n�Ѻ�.F�F�	@���ND�NB�iB�&���|ܥ����o�,3�K���0B6}�a���
�@�P(I)T�%*�J�����|�(�J.�A������������������������kkkkkkkk[[[[[[[Yqqqqqqqrbbbbbbbaqqqqqqqs[[[[[[[Yrci��E*IQ333qqq0w�KF�o"À* %��LA	AԆ�H�ٙ�ِ���,9/B��!Fc��%R���G�H_�Xδcd�����T�	�B���Z4:u:�ӑ��������������������������������D�g&'���&&&&&&&&&%�$��"#��2RW���8�x)���l`���LQ0(���
ƉR�Yr��I(>��E�Q_J��P(<�+��.���3
�����o�������Ԥo_��ڈ"��]�"7���XJ�_};RE)7&�A_�%(�r�R�	}���M��t6�Xt��t�������E)DA�|�7�o$M�|�7Ҕ��a�`h5�a�`h5�a�ph4a�S|�F�D�ݪ�a$���}��p��t7F���B�)B�.F�)B�&��y��ɹa+�A$M����Xw%�pm�v���`�B6�gؠP(
I$��J�R���D�Q(����E��t:�335�����������CƳb��j�jIqqq�����a�	�q�i�I����
�������2.J�(����I'� �+�S�H���"F�`t���D̨z@�7��eJ�*A񙙘��eJ�����:�
'N�h�	Q$ɐT��(N�B�
(P�hM�ө�4X��s��������������2!QRS����󓓒RRRRRRRS��2W������"""}>�DB�c!�CI$�c�I(]
-�+�I%1����B�L����L`0�p\�rXph4�aXw�a�d�~;Qo�j�F�o]��J&���t���nXJ�$�F�i}���Mɺ}� ��
�a+��M��/F�5'U��1�S⋂���B���$�" ��r7W�5�$W���������3a�f��Xv��A�3
o��"H���v��ܛ�BH_}��q�E�^E�]��F���u�M��>�!$)E(��� �)JR��;��8.��`�`�B!�g��(
�@�IJ�R�U��|Q(�]�D��t:�335����������ִƶ������CCCccc�#�b���d�����#b��������E�̒`�6t%K�.K�\,�x�h*� d��
��	cSf*L�%D�*$���bI��zz�UD(P�:u�%J�&LIS�P�:�
(P�B�8��P�d��ҭLOOO�����OO��LK�_B ���g�'%���%��'$d���"#����������22S�2RW�舉�JJ�"1R]b0R�mmm��n/�AE��IQ(R�RK�!v�W�����]� ������$���ȻK������>�Qa�v)��$&�4�48KP l,0م}Ģ��O�ט�Y�T� B���%��w��;��-JO��7��a&�o��BHW�°�y"H��K
°�+
°�04a�`h5�aR�}�JF�j�]��7����R�Q7$�������>��>����}��$&�(������H��K
a�w%�p�v���`�B!>ϳ�P(
�$�IJ�R�����Q(��E��000000qq333333QQQmmkkkkkkkkQkLmt:͍�؍�TM�����������Ϗ����"I�q���%��yJ-H9A���fLU "&AQ!]��bd��� @H�o�I� @���J�fSSf*�
'N�*�
�D�T�ӨP�h�
(P�B�KE�S�N$�3����jjjjf'������&$�� ��g�DO�S�������22222223���2222RW�蔔���D.���}����-n/��``�g�l!�����p�%�p��v��7�$�o��r�u�Y����	�
 pp`c`�I��z8C��,��(����׶Ä9��l"�^b��``p����		z�C�KP	$�t��RBHW�� ��A�D�JR��)aXV�a�f�a����JXv�v��A$R�Av��/��R�QJ)Dܛ�BHI	�7)E�������F�})aXf�r\�y^P`0�F�g��}��$�I$�I)T��|�_J%C���t:\\\\L���TTTTT[[[Z�SI)V�F�c�����cc������c�#�����$F�cdĔ�rch�����(���"1?Wc="= u�QQ�Q��31�J� LH�
�ɓ$�S�J�|cc u
'N�*T�ӧN�:T�ӧP�B�
(P�B���V�έ:��@�����������鉉���y��Jrb*DJFr^JFr^bbzzFFFFFFFF^^bb^^^^FFFFFFrrJFFFF�"%}��" 1:I$B�e���!��g��7ݫ�$A��$���0(*��+:��/QG��`��$8$880�,�z�<Ko0�瘳�9��	x�\������XY��z�;/ ����Q�,4���$)K
�}��
�v��A��D�7Ҕ�)aXV�JXVa�V�������$I�Av��~;Wj���_��/����Do$I})aXf�r\�y]�l�D#a���}��$�I$�R�T��|�(�J%C��`````��ff�fff���ڢ������֘�������h�\fIkIk(���$�� ��*����W"�[e�fj ��?n`(�������3H91cT#WWfHSSHc#c|HT|*L��bJ�fH @�S�N�*TI��eP�:t�R�J�:t�ӧJ�:u
(N�:t�ӧ_��:���L�����������yy���������y�X�蔌�,,U�F^bbFFFFFFFF^^^^^^^^JFFFrr^^FFrrrFJ�}�����:@]/�WA@���y]���a�T��aXV�p
	��jM����s�XX$$8$XX %�,�	z�]��s��4�p��CF��CE��ǫ�P`\Q��		w
<�\/7����,�Rl8^�%�i�S|n��;U�HW��_��ڈ#x�o������,+
o�,+��3�aM�D�JXT�)7�DoD�o�ڻWj �"�7��y"o�)K
�0��k��8.��`�`�B!�ϱ@�P(I$��%*�J����D�Qt:\\L������T[[[[[[Z����ˌ�Z�
�n�cCcCCccc����D���Ud�J������� l����?cH{s1?SB�r�U����P�!\�5E5v3�ٟ٘��&$�5u5vbeN�:t��dT�ӥJ�$IR�N�B��ӧN�:��ӧN�:u����Q\��S�	
��g��g�%��'�f'����'$ddg'%�&'�O��))��������)���y))���y��yy)(8[蔕��}��6w$��e����0��A�h0Y��p�<^�Gc�0Y��z��=^�Qa`�`H����H����  z<\"��7���..�z��oWp��0$$$889�X�z=��������I�E�W�7,%�������ID�7���)JM�}�a���kÃA�3
��)K
¥&�"H��y�H�$��7��	"H�$�"H�$�
°�04ð��༮۶D"��l�>��@�I$�R�T�U|�_J%����000qqq33QQQQQQmmmkkkkkLLL..........4k.Q5w�؍�͊&ɇ��Ɔ������k���Uc���t��$4E�,��UP�����1*���U
�?S�LJ�3�2d�ل�TI3ԅrN�*T���*$�ӢD�&L�1'N�BЩӥN�:��ӧN�:u��!�M��0�-���OT��NNLO��LK�H��ILLO������OLLK�NH�NNNNNNH�D���dg'$��ddde��g%���$d���P001R!QP�p1W�����͸��(�3�8C.�gs�%��		z���盹��					w;��E��W��HHHs��,�,p���"�7s�X801�,,�y�;��7��`  `�c��� x�6�E��G�Ѱ�Aa.�7t��R�	_��~;WjH�$��o��JRH��+�A��kÃXd��aXT�)7��o7��|�$F�o$ID�$ID�a�`h4ð�;��/+�D"�l6}�b�@�I$�R�T�U*�_/�%����0000qq33QQQQQQmmmkkkkkLLL...........Lk.kM}*��1:�͓�����ÛK�|j�	D"x�Ul+�����)��*��̨U��	�����f5vfff4����i
o�ٙ�	&$��	*lo�N�*$�2ʕ:$�ҥD�&L�1%N�hЩӧN�:��ӧN�:u����Q\J��T�����LK��O�LK��OO�K�NIIK�O�����OOLLLK���N_O�RR23����23��3��2222RRRW������XXX888˼\9�4X �, 	z��n�s���w;��W���,,,,�z�^�W����p�\!�"�Ws�P]��w;��W����z���8@ /����x�9UD.��Giy�7)E(�����%��	�a��a\l�0�3
¥)K
°�+
°�+
°�+
°�+
���"o�,+ð�K����n�0!�D#a���}�g��(
�I%|�_J.�C���`f��t�����������������8��6��8���(�]OC̞�'���)�A��_=�&���5���EIK�O�K�T���ٙ���ٙ����f| L�2�3+��&���LI2J�&�ƨ~���LIS�P�:t��(N�:t�R�N�:t�ӧP�hѡӥI�h�:o����Ϗ��
�*u���!!!QQML���ļ�����������䔔������������ļ���䔔��������ļ䌔��������䔔��DD**DDDDD****2�z�K����!!������		z�^�Qaag����z�^�W�HHHHHpHppppp``c�8$Y��y�
;�����,,�z�����8\.����z)9^�Oh�����ȯ�~+�ܰ�E�$W��A�)�H�A�3�0�+
°�+
°�+
°�+
°�+
�0�I�o�,+ð�;����n۶D"�l6}�g��}�I$�I_/�%����0qq3Qt:L��TT[[[Z�������ˍ��[Z�����O��LNKIB"�F����� ±��]���
%S%1SHcWcTSTTHHcccccWf|||ff||fff|&M��2dɐ|| A�]]�I7�g�"D�*TI2
�
o��	�*t�(P�B�
'N�*T�ӧN�:t��4Bt����B$����	�:t�666664��E53���3����3����茼�����������ļ����䌔��DDFr^^^r�}��������DDDB�DDDDDDDDB���aa`b��c  A�@`HHpHs�XXXXXX$$XXXXXXXXXXXXXXX$$$$$$$$XX$$$8888$$Y��y�����XXXXXX$$$8881��p�   =����CCM��a��l6%�Q���1��x�<���r�&���K�ݪ�J,%ڍ��R����h4a�f�A��h5�a�f�a�fa�V��Xv�r\��p�m�v����B!�ϳ��
�$��J��%����t������������������������6��5��5�16�[]ͦa�CLAL	�Ź�DuSw�����+�$1�33+�*1������3+�>> A�����2dɓ&L��3�o���� �@IQ$
�*$��ĕ*t�(P�B�
'N�*T�(P�B�F�4ht�S��BT�2dĉ*T�-+��������*)��������O��H�G%��dDD�&&'�����秦&&%�����$o�!QPA�R3��2PA2"2222RRRW����""""""}>���EEEB���Ȉ�FB��BC� ��!"��W�HHHHHHHHHHHHHHHHHHHHHHHK��,,,,,�z�^�Qaa`�����������  ����z;��Õ��r�\�W)c�����Z�x����Q��l"���گ��H��%���� �,;��0�04�Xv�a�v�a�f�a�f�a���0���r\�%�p�vݷm�"�l6>ϳ�P(	$��U*Q(�]�A�������E������������������\�QA6L4>4mLQLqqR@O��WΑf|�U�ږ��B_��ULU�$1��������33333>>&L�2o�����	�*T��d��A���Q$	*$���J�&��LH��N�:ѣF�4h�
�N�*�
(P�BѣD�!:��t�Н*T�ӧP�B�:u������lli	
�jg积���53ӗ��yy(�Y)yy���������鉉yyyyy�+�T(���*"*DDD�}>�O����***DDD�%"""
w8F��G��08$$0888888888888888$$$$$$$%��z�����������8\  G���XXX4�v6W+��ZZZZZZZZ�r�[-�+a��l��"(�&����҅�^E�D�o$M���aXV�a����a�v�a�v��A��h4r\�aܗ%�r\�p\�vݷl�D"��l�>ϱ@�I$�R�U�D��t:]
*.����kkk[[[[[[[[[[ZaE1�ͬ����fQ.^"np�� ��'q���\�[&ΕE2���eC�����F5F64��E3��fffg������bD�&L����D�*t����ĉ&��L���
�*LH��N�L�R�N�:u�F�4hѣD(P�:u�F�4hѢu�V�Bu:t�ӴBu
-4N�jիU����������K�T��K�NK�IB��_G'%�'�����秧�&&&%���$dd���DAc ��"!���# �`aaab���`ab�DO�����XXX��8X��8{�4Q��x�@  .���p�\.�������������������,,�p�@  /�����c���r�[-��iiIIIIIIIJ"�k���r�[���aJ�K��7�Dn��B�����W�o�,+��;ð�;ð�;ð�;ð��ÃA�;��9.��8.��n۶���B6�g��$�I)T�U|�t:��k��Y�������֘��������\�\�Pq4(:\\'���%�xZ2�µ����$gꏌ�'�i�'�
ꇯ�����������Ϗ�����ĉL�$H��J� �$�Q$	:$�eJ�LIT(P�:�
�N�:ѣF�4hѣD(P�:�:t�ӧN�:իS�B�:t�4hѣD�ӧN�jլlli		
��li	
�jg秧������%�/��p1R23������������������2 ���B 0GK��
"""22DDD*D*22"22".�	 x�\.   ���p���������������    <^/G��ӱ��l6��d������III흹��)ggr�<ܫ���sPi��	���F�D�JXV�A��h4a�v�a�v�r\�aܗ%�p�p^W��vݷl�D"��l�>ϱ$��J�W�����000qqQJ�����������&5����������A�
Jɮ��;���Dt �Q��FrD��Fb��~b�Ʀ~���ƮA�����2l��Ϗ��>&LI2dɓ @�1%I�*T�Q$ĕ*$��J� L�ҢI�:��F�4B�
�S�N�:t��4h�
�S�N�:t�ӭZ�jv�V,Z��t��4h�:իS�Z��!!!QQQQ]�!!QQMMML����ML���*FFr^b~~~~~~zzzbb^^^bbzzzb^F�"""}���BHP((���8X�XX888�88XXX����Ȉx(8xP�9�        �p�8\!��!!!!!!!"��!!!���!�����pppp``c� ��x��Gc���l6�R���Ғ�%$DDDDDDDG4DDG7�Vw7Vw���K���`i��z=\F�tn��R ��y����04�A��h5�r\�%�r\�%�a���h5�r\�p\�y]�m�v����B!�ϳ��I)T�U|�_:�2J�[�[Skkkk[Zbbc[[[[[[[Y��i@l�,��x(D^�2�z���|11W|9 z~��$�3��B����euuvbĳ333>>>| L�2dɓ&@�eJ�&$�ӥJ�*T�2eN�&@�S�D�u�F�4hѢ'N�N�:t�ӧhѢ(N�Z�jիV�Z�b���X�;D�V�h�:t�V�N�j���BBB����������������A��)��Xz�A��������鉉y�)��������XXX#�P\ <,D<��
"
t����O@  �����008$$$%��y����8\. ����x�^/���XX444�r�[%������*JH�noon������N��Ψ�mL*���ML��ҕ'��+���|�/�7M�"�W�°���R�"��;���+��K�r^Wm�a�w%����6�l(��a���6pXW �P�A��$�I<����Q(������Y�Y@�l������J�������^**�t�����LOU��LOO����و�������A���dɓ&@�	�&LH�%J�*T�R�N�:t�ӧP�B�
(P�B�
(Z4h�:t�S�N�:t�ӧN�:t�֭Z�jիV�Z�jիS�Z�bŋ�Z�jիV�X�c&L�,X�]]]���!!QQQQQQQQMMMMMMMM�PČ����D**�9?T??SS??=1?111//9999999999}>�B���EB�AB���C�]! @0�@@�K��2"2""22�t�;��/�```ppHHH��HHHH��$$88000001��p�  <^/����x�;��+e��----))RRDss{uugggjjjsj``gugM`)^nnPsouD{u{jjRDr�;��A�����޿��"o���ÃXbE��)JR°��R��K
o��;��r^P`1�^Pc�6%J �������B����&�AE|�It%J	W����$��r�]W[ܡAB���/��y�,T��ļ���QQP����MMQ!!MQ!����uuuvg� L�d� @��dɉ$�S�N�:t�ӧN�:t��(P�B�
(P�B�
�'N�j��ӧN�:t�ӧN�:u�V�Z�jիV�Z�jիV�X�būV�Z�jիV,Xɓ%�,WWWWcccHTTTTTTTTSSSSSSSSccH?/#9/9#}>�NOO�O����LK���OLK�NNNNNNNNNH�H�EEH��D@c!�# �" ����Q�WK�`Q�2"""2
�t�����  .���HH`````p``c���p�\   �İ���������v6�+���l������)"9�����555777&�&��&��.�=�0(%�7���3���7(9����(�y7_|AJ!}��nW��XRD�aI)p	�7���J]��v��(8 ��(0�� 1*�Qy\ؠ�7�A���B��v�i�����'�0" �'s��č�Jrbbbbbz~�b^^z���zzz~~�������Ʈ���������@�	� L�1$ɓ @�2dĉ*T�R�N�:t�(P�B�
(P�B�
(P�B�F��Z�jt�ӧN�:իV�Z�jիV�Z�jիV�Z�jիV,XɒիV�Z�jՋ2d�vL�2ffWWWcccSSSSSSSSSSSSSSSSHcWT/}�����������������������������������������DDDB��``aa`��N��@��!qGK��""2�x;�N��'���z8@/G��� �   x�^/����z6��a��l9\�V�d��������III���՝����555���yuuAAAA�-Y��u�5y�%�--��y�t�-���|fI$���	��0��$&�a����}�B����9.H��Xg$BI}�W�p�H4���W r\���}��m�}��m�-y�9&j�j�ƍ��A���ҙy)�;茼���T�������ļ��Q!L����MQ!!!Q!Q�]�������&L�2dĉ&L�ĉT�R�J�:t�ӨP�B�
-4hѣF�4hѣF��N�jթӧN�:t�V�Z�jի,X�bŋ,X�bŋV�X��&K,X�bŋ,dɐ�dɓ332���������������������A{蔼���ļ�������������䌔���999999999#%}>��@�adDDDDO��x �888�x (S�44 (()��t���@A�DC����PP@h����x�;��`h���z;���a��l�[-��e�ZRRR�����������������ܚ����������ޠ�ެj�j��j��������pj�pddx�p��j�� 8EgUVjkA6$�+�D��}�ϳ��Xw)$Xw�7�m�p]�m�p] �
��$�j.K�IpXW%�a�K��d�R"*��Z��p��@�DAEA��LLNIIIE@���H���T��D�&&&'$g�&'�j��g�j�lj�ilj�Ϗ����&L�2dɓ&$H�"I�&LH�%J�:u
(P�B�
(P�B��F�4hѣF�4h�:t�V�X�jիV�Z�jիV�Z�bŋ,X�bŋ,X�bŌ�2u�,X�bŋ2q�dɓ'�ffeuuuu5555555555555553�F4���������������������2W���rrrrrrrrrFJ�"""}����>�DO�R 0p1P00000ppp�xk��
�w;�B�]!@ ���  !A�xh����w�<Ń���+���l;��a��l�\���d����������������������՝����55�yyuAAA�-AT���T�T�X�ѭ,����\�����j��7:�����YފHa�M��z�驙�U�}�t ��
7��3��iH��J���l�\�H�`�m�1E�6x�=FAȝ������$�/�#��y�x�Y�蔔���D*rzz~zr~z^bz~�~zz~z~���Ʀ���Ʈ���̮����@���	�&L�1"D�$H�"I�&$IR�N�:�
(P�BѣF�4hѣF�4hѣF�4h�:իV,X�jիV�Z�bŋ,X�bŋ,X�bŋ,X�c&L�u�,X�b�L�8�ߎ8�>333+�������������������)�1�������������������������������������������DDB�b�DO�1R" �0� ��00pq�����)�((.�t����K���w��@��n���i��------))RR)RRRDDDsDDDDDDDDs{{{uuugggjjjnnnnMM`^]]PEEEoooKK8UPEVIAb@.I48g@2m,D4E{V26Vjv7��<�n�GӕY��)K
	l6���(%��l%�k}���(�	H1�NV��I$̢�6�B ���w�x��dU�J�"=%1S#}>�LO��H�H��ONH��K��������|||| L�7��	�&L�1"D�$�R�D�&LIR�N�:�
(P�B��F�4h�:t�ӧN�:t�ӧN�:իV,X�jիV�Z�bŋ,X��&L�2dɓ&L�2d�b�L�q�2dɓ&L�2d8�߿q�|||ffWWW????????SSSSSSSSHTSc| ��^b~����������~~z�~~zbbb^rrrrrrrrFJ�"}���B�ȟB b�``ab�a``�!��" �  ��!@�O�� PP\`5��x<�b��K���w<�o1AA��K��Z��R���������������������������������ܚ���������������ޖ���d���j�x��`|h� ���j^#
w��F ���# /1g)����z�W��W���I$n��fq��v��^��*���,��D


t�� ����������������1��������������$*)�$1��**1�fcccW| L�2dɐ&L�7�&LI1"D�*TIR�J�$�R�J�:�D-4hѣF�4hѢt�ӧN�:t�ӧN�:իV�X�bŋ,X�bŋ,X�c&L�2dɓ&L�2dɒ�L�8��2dɓ&L�2q߿~8�TK�BC����ĽP�����BBB���C3�������yɉ�������y�����yy��)))�y興���,�T��d�,<<d,TTT,DDDD<d(\!�.�x;����  � �@�x����1�(�w���XY�Y��/onl���on������
Oi�n����mJ����J����/i*�OGC�8s;�c��)x�
�������������������:B��CB.�q@'��`a�,�w���Wp���h�g>.x<Ɲ��K���t�@@A����DFA��H�Ab��3����������������EEEEEEEF665uuvfb @�	�&L�2dɓ&L�R�J�*T�R�J�*T�R�J�*T�ӧP�BѣF�4hѢt�ӧN�:t�ӧN�:v�P�B�:իV�Z�jŋ,X�c&L�2dɐ�8�;&L�2dɓ&L�2dɓ&L�2dɓ��߿~���9�$���ُOT�NO�1�����1���3>>>3������������������)��������������������������D@��A�@�I_B�`a`��"""## �  #.���H���x��C^ �/�@ !Ap�H@��$0%�,� z6Qڙ�[����[����XW[�W��WTQWX�WXڐ׍W�R��]��nP�F��8��!�p.�-}
����������������� �:]!A@N��h��C�`Q�(0�x;����/ �Q@PЧK���
""}����������������������$$$$$$$1�����33 @�&L�2dɓ&L�2dɕ*T�R�J�:t�ӧN�:t�ӧN�:u
-4hѣF�'N�:t�ӧN�:t�ӧN�
�ӬX�bŋ,X�bŋ2dɓ&L�8�8�dɓ&L�2dɓ&L�2dɓ&L�?~����ߎ8�:M�]������P����x���2���C1j�	i
�g�
g/��zC2��B���yɉ�����y��y����*�##=1
w��;�Awx�@xk��U��z�����ޯWs��,� v"50(/)"7��5"�0&��(7����7��0%���������1*�+6[ �V'�H��XY�`�XA�(Xx( XȈxxx�Ȉ S���x;��B���с�ч���!��x:^ ��P�Wx @P�((((DdDDdddTTTTTTTU�Jrbbz~z~~~z~������������������Ʈ�������@� L�2dɓ&$H�"D�T�R�J�*t�ӧN�:t�ӧN�:t�(Z4hѣF�4h�:t�ӧN�jիV�Z�;D(Z'Z�bŋ,Xɓ&L�2dɓ&L�2d8�8�ɓ&L�2dɓ&L�2dɓ&L�2d����߿~8㎝�Ro�	�*$�Us�%_��K�����ff|||fcHcT=11ScfcW|&$�2i	
�������������1����������������>�@�H�B�@Ȁ��@�@��A�!AC N�p��k���]��x=E	NEb���w��a��v�5;]�M�
���˪���jJ�
�

Ʃf���gǉe�i��!�7ӱ��rzbD�//9}>�FINK�H�C��EB��DDDDFD@]!���xhh����h��4Pa�0(..(..�y��E�@��H(((x8X88XXXY)))+��DDFrb~~�~~�����������Ʈ����Ʈ������������@�2dɓ&L�2dɓ$�R�J�*T�ӧN�:t�ӧN�:t�ӧN�:t�(Z4h�:t�ӧN�:t�ӧN�jիV�Z�jv�4N�bŋ,X��&L�2d�q�q�q�q��&L�2dɓ&L�2dɓ!�q�~����߿q�X�	RbJ�$�,�V�*M�]]��t�7¨I�TI2�j�ό���ĕ:t�����ςN�HS??ST?1=1W|?99}*f1"91"9=/"%=1#x����]!N���e�L	�JD"�
"=?
y�<ޢ�!GHS�%��#x�9�7�������(.��($�����%���L�-I���lj�$jj���b�b��P�Wщ����,U�D*22�w���@�CCCC@�^�q��h������81��
t�:@A ����A�Ȉ��EH����G'''$dd��%��j���
��ilj������������������Ϗ��&L�2dɓ&$H�"D�:t�ӧN�:t�ӧN�B�
(P�B�
(P�B�F�ӧN�:t�ӧZ�j��ӧZ�jիV�Z�;F�֭dɓ&L�2dɓ&L�2q�q�q�q�dɓ&L�2dɓ&L�2d�q�q߿~�����q�X�	R�P��:-�h�;D%D�*M��J�P�h��R��N�:M�D�S�h�����'Z@�2d�	�T=?%99/WM�ļ�]P�Q]�!��L��~DDJ*�}�WffH99TWc1y�  ;�^���G���c�P��( R�n^oV@5KoKbz��� ���*�3� (��<ޯ32��C�23�5E3�2"7��LĈ��JFJ�}�����B�����C�B�.�HP@C���w���B��{���w�;Ȃ��DA@�B��Ȁ�����_D�O�RRRR23����������5EEED��D��65vfffffffffg���������	�&L�2dɓ&$H�%J�*t�ӧN�:t�ӧN�:�
(P�B�
(P�B�F�ӧN�jիV�Z�jթӧN�jիV�Z�jv��Xɓ&L�2d8�8�8�8�8�8�ɓ&L�2dɓ&L�2dɐ�8�~����ߎ8�d��-�:�kB�ѧZ�būS�ht�S��Z�bt��:Ѣt�2dɒ��N�BTH��Z'B�
'J� T����ʛ31���0��Y�>>&$��ٙ���SScTTS/fT�AS�_�f r�y���C����K31(;��� r��� *����*�"�1"��$�5"��A@C��T����ONORٕNO��O�LOLINK�IH�ONNI_DDDDDB�`�#### .�H ���
x
;���B��A]!P!p�QQ 0�P��8)興����������似�����������MQQ!!!�!!!��]���������� @�ɓ&L��"D�T�R�J�*t�ӨP�B�
(P�B�
(P�B�
(P�BѣF�ӭZ�jիV�Z�jիV�Z�bŋ,X�jt�ӭXɓ&L�2d8�8�����߿~8�8�ɓ&L�2d8�8�8�߿~����߿~���:1�'h�:֍�h%�5�V-d��$��4h�:u�2d�:u�S�Z���߿bt%_��;D�V-huF�J�*��B�2��A4'X��U��BU�!��2d	�BLK16�Uʴ||LI�3(U�ʉ|:tI1$��������1���E�HT#y�F"���V��U`B��;{{:����xQ��P���L����PĽ�!!!QL�����L��L��ļ�����䌕��}�������O���P��PP�GH��P<��
x;ޠ�/ w�Y)��x�<�䔕��}���������������$*�����$$1�$*$1���3333333&L�2dɐ @�2dɓ&$H�"D�*T�R�J�:t�(P�B�
(P�hѣF�4hѣF�4h�:t�V�Z�jիV�Z�jŋ,X�bŋ,X�:u�8�8�8�8�~����ߎ8�8�dɓ&L�8�8�;��߿~����߿~8��vK�d�vKZ4Z�w����~ɒūV2vL�,X��&L�8�8�߿dɓ&L�2Z�jթӧh���$�W|TIuF2Z!*$J(P�B�	ӧN�:�	ӧJ�*$H�%J�*T�(N�*TI2d|||c �zr~b*"@���y`pXS�¼�Ίl���Rbz�C�H�FFT��X������������O�OOLLLLK�NNNH�D��d��!P0q����@@@@�����@@�P�2"R22RW�蔔��似���ļ���������MMQQQQ!!QQQMM���]]]����������&L�2dɓ&T�R�J�*T�R�J�*T�ӨP�B�F�P�h�j(P�B�
(P�B�
t�ӧN�:իV�Z�jիV�Z�jŋ,X�bՋ2d�q�q�q�q�w�߿~����߿vL�2dɓ&L�q�q����߿q߿F�4hѿ~;%��2~�bt�?~����߿~;%�V�d8�2X�`�q��!�w��2dɓ&L�,X�jt�Ӵht��d�	�:t�7��)ִ*$J(P�B�
(P�B�
(N�*T�ҧN�:t�ӧN�:t�$ɓ&L�3�����Kɳ$	}8^#" `Oi�mH��� �/� wл`%��HH}>�ɤ)�1��**$1�������$$$****)�����������������������������DDDFFFFFA��������DC��AB�Dg''$d���)�yɉy��������������������BBB�������333333�� L�2dɓ&L���J�*T�R�N�:t�ӧN�B�
(Z4B�D�P�B�
(P�B�
(S�N�:t�֭Z�jիV�Z�jիV,X�bŋ�X��&C�8�8�8�8�~����߿~���dɓ&L�2d8�8�8�߿~�����4hѣF����ɓ'�X���߿~����ߎ�bի8�2X�q�q�q�q��&L�2d�bŋV�N�jt��%�֍!:U�խ
��
(P�B�
(P�B�
'N�*t�ӧN�:t��(Z4hT�R�D�*u�v7�τ�OΤ����K[��*��s� �j�ll����ɕfc ̮���Ʈ̮�����ƐƐ���������~~zzzzbbb^^^^r^^b^rFJ222***DDD�}
������������������������������������������*$$$1���$$**+����3>>>>>> @�dɉ$H�"D�*t�R�J�*T�ҧN�:t�(P�B�F�P�h�kF�4hѣF�4hѢիV�Z�jիV�Z�jիV�Z�jŋ,X�bՋ2d�q�q�q�q�w�߿~����߿vL�2dɓ&L�q�q����߿q߿F�4hѿ~����2~�q����߿~����X�j�O�vL�,q�q�q�2dɓ&L�,Xɓ&K-Z�jŉӡ:T�1�Z'N�:�KU�F�4hѣF�4hѣD(P�:t�ӧN�:t�ӨZ4N��ӧJ�*T�RiϏ�Oо���>)��� ��>1�TW|SHhu� K��S����>3333>>333+���������$****)����������������������
��������O��)))���""#/1=1==1//1======?=????SSSSSSTTTHHHccWcWccHHHWfff|||||| @�2dɓ$IR�D�*T�ӧN�:t�ӧN�:t�ӧZ4hѣF�4B�D�Z4hѣF�4hѣF��Z�jիV�Z�jիV�Z�jիV,X�bŋ�X��&C�8�8�8�8�~����߿~���d8�8�8�8�8�߿~�����4hѣF���ѿ���ߣF����߿~����X�j�O߿vL�8�8�8�,X��&L�2dɓ&K,Z�bթ�!:U]��S��Z�vM�BѣF�4hѣF�4hѣF�P�:�
(P�Bt��(P�h�	ӨP�:T��2��1�3�Bo�$g���AB�i�2j�Ī31��&��L�2�_� A���o�����������lli			
��jjjg��秧�&'�����%䯢!P��R'����%%##9##%}
������������������������**)�****$$$1����3+������3>>> @�dɉ$H�%J�:t�S�N�:t�ӧN�:u
(P�B��F�4hѣD(P�Z�:t�ӧN�:t�ӧN�jիV�Z�jիV�Z�jիV�Z�bŋ,X�jŋ2d8�8�8�8�;��߿~����ߎ;&C�8�8�8�8�����ߎ8�ߣF�4hֲ~��%��7�~����߿~;%�V�d����ɐ�8�;��d�j��2dɓ&C�d�bŋV�Z��ӥY��	�B�:�L�4:��F�4hѣF�4hѢt�4B�
(P�B�
'N�*T�ҧN�*T��dēWc|THHcWfffc��%��<�1�U�г&L��1/�ʉ&��@�2��	� A��񙙙���]]���!!QQQQQMMML���������L��Č��DDD�}>�D���dde�'$d�����Fbz~~~�~zzzz~�~~�����������������Ʈ������̮������@�2dɓ&$IR�J�*t��(N�:t�(N�:t�ӧP�B�
(Z4hѣF�4B�E�S�N�:t�ӧN�:t�֭Z�bŋ�Z�jիV�Z�jիV,X�bŋ�X��&C�8�8�8�8�~����߿~���d8�8�8�8��w�߿~�q�~�4hѣF�h�߲Nuc'�ѿd����߿~���-Z��4oߎ8�q�q߿�ũ�2dɓ&L�;&L�-Z�jv�N�@�1%N�N�j��P�Z�:t�ӧN�:t�ӧN�:v��B�
(P�B�	ҢH>>*t�R�J�f|:MP����BC3��A�iI��3Ubr�I�L�Ӫ�P�&LH�d>>&L�������������������O������LNNI_O��))���yyyyy��+���%91=???S?====?SSSSTTTHHHHHHHHcccccWWWff|||fffWW @�dɓ&$H��J�*T��(P�:t��(Z4B�
(P�B�
(P�N�:t�ӧh�
-�N�:t�ӧN�:t�ӧZ�jՋ,Z�jիV�Z�jիV�X�bŋ,Z�b�L�8�8�8�8�����߿~����ɓ��߿~���8�;�߿~������hѣF�쟎��U���F����߿~����X�j�Hѿ~�q�8�8�~;%��4dɓ&L�2�&L��Z�jv�J�T���Z'Z��v�P�d�:t�ӧN�:t�ӧN�:v�!B�F�4B�	Ҥٕ�ʕ$H�"U��	���' ������~��ev�	ʘ�f ��]�ӯ�eZ&T��d�>>&L�2>>>>>333+�������$****)�������������������IH����LOOOK��NH�I_O�S�����3����555EED��D�4�4�66665uuvffb�������&L�2bD�*T�ӧN�B�F�N�BѣF�P�B�
-4hѣF��'h�:t�!B��թӧN�:t�ӧN�:t�V�Z�bŋV�Z�jիV�Z�jի,X�bŋV,Xɓ!�q�q�q�q߿~����߿~�q�2~����߿q�q�~����߿q߿F�4hѲZ�:�L�-X���ѣ~���ɓ��ɓ&L�2w�ߣ~�4hюɓ%�,h�`�߿~8�d�bũӡ:$�"J�*t��K-Z�;F�4hѣD-4h��T(P�:t�T(Z4N�j�%J� ̮�L����ʇ����dd>>33+��&L�bD�*T�S�N�:t�ӧN�B��ӥJ�$�2d&A�����������]��!QP����MMMP������������䌌�����������似��ļ�������QQQQQQQQMMMQQ!!!�����]]]����]]]]�� @� $IR�N�:�F��N�:t�ӧN�
'N�*��v�ӧN�:t�ӧN��ӭ�N�:t�ӧN�jիV�Z�jիV�Z�bՋV�Z�:t�ӧNѢt�֭Z8�8㎱bŋ,X�bŋ,X�jիV�Z�bŌ�2d����߿~�4hѣF�4o߿��-h�c&L�,d�w��ѿ~�q�~���ɓ!�����q�q�vL�,X�:�߿~�q�2d�būS�BTI4�ӧZ�jիS�B��իV�Z�jv�֭N�
�V�N��A"J�:�D%J� ���t�ӧJ�*̐���L��33�ĕ&L�	�T�R�J�:T�R�J�:t�R�J�*TH�$ɐ&@��32��33333332���B�������B�BB������������鉉�yyyy��������yyy���������BBBBBB������BC33333331��g�ffg��������dɓ&L�2bD�*T�ӧN�B��D(P�B�
��Bt���ӧN�:t�ӧN�:t��h�jt�ӧN�:u�V�Z�jիV�Z�jՋ,Z�ju�V�Z�j��ӭZ�b�L�2dɓ%�,X�bŋ,X�bŋ,X�bŋ2d�q߿~����ѣF�4hѣF�������'N�q�2w�ѣ�F����F����8����h�q�q߿~8�d�j�߿~;��vL�,X�;D'N�X�c&L�ɓ%��Z�jիV�N�jt��!Z�:t�ӴhѢt�ӧN���D�ff||| @����g�dɐ @�"I� LH��J�:t�ҥJ�*T�S�N�*TH��J�L�2���ٙ������������������OOOLLLLLLLLNNK��LLLT������������� @����������ɓ&L��$ĉT�R�J�:t�'N�:t�ө�4h�
)ӧN�:t�4hѣF��:�:��V�Z�jիV�Z�jիV�Z�jի,Z�jt�,X�bŋV�X�c&L�2dɓ&K,X�bŋ,X�bŌ�2dɓ&L�2d8�q�q�F�4hѣF���:4hѣF�4hю�:�Oߎ8�߿F�4hѣ~��4h߿~8�8�ߣF����߿~����u�Y�q�?~8�d�u�-NѢt�ӭZ�`�d�bխ4hѣF�P�h�	R��4h�
�4h�:t��:TI2eJ�:�
-
�WcW| @� T�Q"J�:t�ӨP�Bt�ӧN�:t�ӧN�*t�R�D�&L�2���Ϗ������������i	����jjjj���������秧�&&*jg����秧�����jj���		llllllli			llj��� @�ɓ&@�ɓ&L�2bD�$IR�J�:t�%N�:�
(P�B�
)Ӵh�
)ӧN�:t�4hѣF�Е:�:��V�Z�jիV�Z�jիV�Z�jի-Z�:t�,X�bŋV,Xɓ&L�2dɓ&K,X�bŋ,X�bŃ�8�8�2q߿q�q�~����߿F����w�߿~����߿~�j�Oߎ����ѣF�4oߎ:4oߎ8�d�q�~�4hѣF�7�ߎ8�V2q�2~�q�dɐ�d�jթӧN�jիS�h��ҫV�Z�jըZ'N�	ҭ4h�
"D�&L�2bD�&@����%J�:t����C����Z':��R�P�B�F�ӧhѣF�4N��F�P�*T�Q"I�*TH�d @�&M��]]MMQQ!!!!!!!!!!!!QQQMML���!!QQMMMMMQQQ!!QQQQQQQ!!�!����!!!!���]]]��������2d @�2dɓ&L�2dɓ&L�S�N�B�
(P�BѣF�4hѣF��Bu�F�4hѣF�4hѢ�Z4N�jիV�Z�jիV�Z�jիV�Z�jիS�N�bŋ,X�jիY2d�bŋ,X�bŋ,X�bŋ,X�q�q�c&L�q�q�q߿~����߿~8�d����߿~�����-Z;��8�8�~�q�d����dɓ%�,dɓ$hѣF�7�q�2X�q�����vL�2d�bŋ�Z�jŋ2d�būS�Z�jի�h�:t��hѣD(N�B��ӧJ�NѣD(P�$�2d3&$�2�D�L�2�*T�S�P�B�F��B�
(Z!h�
'D�L�2
�$� @�|fWWccWWWWWWffWWWWWWWWWWWcccHHcHHTS??=SSSTTTHTSSSSTTTTHcccHHHHHHHHcccWWWWWWWWW @����31 @� @�1%J�:t�ӧP�B�F�4hѢ(P�:T�(P�B�
(P�B�C�J�h��t�ӧN�:իV�Z�jիV�Z�jիS�hѢŋ,X�bիV�Xɒŋ,X�bŋ,X�bŋ,X�c&L�2dɒի2dɓ&L�2dɐ�8�;��;&L�q�q�q߲Z�w���&L�,X8�2X�c&L�,X�jt�֭Z�c&L�2dɓ&L�2X�k%��2X�k��;&L�,X�bŋ4h�:u�Y2d�bթ�4hѣF�
�:t�Q$ĉ&L��:t�Q"N�:T�R�Z:T�2�J�fSSf&������~~$I2	�*LH�%J�*T�R�J�*t�R�D�L�2 A�]]]]]]]]]��!!QML�QQQQ!!!!QQQQQQQQQQQMML��ML��ļ���������������L�QQQQQQQQQQQQ!!��QQQQQQQQ���]]�����������]]]]]]]]�����dɓ&$IR�J�*T�R�N�:T�Q"J�*T�R�P�B�
(ZUD�4hѣF��Z�jիV�Z�jիV�N�;F��Z�jիS�N�jիV,X�bŋ,X�bŋ,X�bŋ,X�bŋ�Z�jŋ2dɓ&L�q�qߎ8�2Xɓ&L�2dɓ&O�-Z�w�X�jūV�X�jիV�Z�jթӴh�:t�V�Z�jիV�X�bիV�dɓ%�V�8�X�b���Z�h�%J�:t���euv67��������65uuv4�EEEE553��EE3�������}>�O�q�������n`u-y�:DITو>>3+��>>33>>> @� @�2d|| @����33��2�BBBBBBBBBB�����yyyyyy�������)))��y�+興����似���������QQQQMMQQMMMQQ!!!MMMMMMMM]���!!!!MMMMMMMM��������!!���]]]������ @�J�*$I2eJ�*T�R�P�B�
-���D(P�B�
+V�Z�jիV�Z�jիS�NѣF�ӧN�:t�'N�jիV�Z�jի,X�bŋ,X�bŋV�Z�jխ'N�jլ�2dɓ&C�8�8�8�,Xɓ&L�2dɓ&IQ�HN�;F�4hѢ(P�B�
v��*$�Q"I�||fHWfcS11=9/1119%}�����A䢢 ���䧧�b��G��j�g�j��$@��� �b���ac!o���R ������K���w����������t�].�K���	,p��BF_F*�lllllllllllj���������llli			
���g�&'�jf$jg�/�QR""22222222�󓓒2223��7�����L�,���� �<-����}>�@`��a���b�O�RR�P2�w��3��5D�vfd��F6g��d���C��555D�65ut$�U�R���������������� @��$H�"J�*T�R�N�:�
��h�:t�֭Z�jիS�N�:t�ӧN�:t�֭Z�jթ�4Bt���N�:t�ӧN�:t�֭Z�jիV,X�bŋ�T9"}��u��Oѿ~����߿~����ߣF�4hѣF�2bV-B��R�J�*T�ӧN�:t꺻B����))+興TT�J*"�/S/% UV)"}�������Li
i
�����jf$o�S��EEE3�S��EC�����󓔄�E53���ffg����
��������j��
�'���j��Ϗ������&L��/��������||fff&�ƨ����A�]P��MQQQQQQQQQML�����􈌼��JFFJJr^J�}����# �B#�������x;��'�)�y���A��*�Euvfg�>31��|W|| @����&$I�1$ɓ*L�2dɉ$H�"D�t�ӧN�:T�R�J�*T�R�J�*T�R�J�*t��(P�h�F�ӧN�jիV�Z�:t�ӧN�:t�ӧN�:t�ӧN�jիV�X�jիV�Z�jիV�Z�jիV�Z�bŋ,X�9W�g�'Z4Z�w��߿~����߿~����ѣF�4hѣF�MM�B�J�*T�R�J�$H�"D�>33+��$ ����̮z�@I2	�3+���*�@�V�
����Z��61(S�ht��o�ςD� $I7�t�E2�$H�5w����|ffL�2WWWWWWWW&L�2dɓScfWcHHc&L���2���������2dĉ*T� ��L�2 M�P�M!]\��B����������������鉉�)y��y��y(XYy)�����d�<`�M��L���y�����\�5s�UEEEEE552�������lτ	�&�����@�	�:u
�P�B�
(P�B�
�ӧN�:v�4hѣC�N�:t��(P�B�
�P�BѣD(Z4N�:u�V�Z�jիV�Z�jիV�Z�j��ӧN�:u�V�Z�c%�V�Z�jիV�Z�jՋ,X�b�L�2dɓ&L�,d;�c���4h�߿~����߿~����ѣF�4hѣF�ubs�
�:t�ӧN�$H�"D�:t�R�J�&L�2d!*�~^~�u	�$ġZ�jr���;FC�h�kA'N�:TI1"I�*t���N�$�2bJ�:T蒢J�*M�bD� A���������2 A����������3����2�3�ɫ��������&L�2dĕTH�dɓ&L����
�o�ɐ||fcHHHTHHHHHHHHccHHHTTSSSS?1=Tcf ���A�L���\P�\���] ��BA+�!��!��]]����)zB��333�
��WH|:��@��"D�&L�2dɴ?S:u\�S�N�:T�ӧN�:u�F�4hѣF�4hѣF�4hѣF�4h��(Z4h�
��N�jիV�Z�jիV�Z�jիV�Z��F�4h�	ҥJ�:�bŋ,X�bŋ,X��&L�2dɓ&L�2d�:�C�~�����߿~����߿~����ߣF�4hѣF�u��&�`��J�*T�R�J�*T�R�D�$H� @��X�A�#"��j�j��P�B�:v����|ft�ӥN�:$�Q$ĝ:t�ӧN�B�	1%N�:T�D'N�*L�bJ�L��"D�T�ӧJ�*TI2dɓ&L�lʊj�
�j�
��ffffffff$IR�N�:t�R�J�*$I1$ɓ*T��I��$�2	�&L�2dɓ&@����BA��)zC�ʢ�Z�)��sB�ȉ(8Ȩ#�(d)��w��o7�����+����OO���S1}3)��$$*)��$$$$$$$>���T*T�R�J�*T�R�J�B�
(P�B�
(P�N�:t�ӧN�:t�ӧB�F��B��D�ӧZ�jիV�Z�jիV�Z�jիV�N�:t�ӧ*TI2bJ�dɓ&L�2dɓ&L�2q�q�q�q�Z�w��X�7�ɒ��߿~����߿~���hѣF�4hѣh"%iR�	�&L�2dСB�
(N�:t�ӧS�N�jŋ�Z�K����B�b�S�����bҬl��N�jօD�t��'N�B�
%N�hѣD-!:t�ӧN�h�	ӧN�B��F�D� ����T�R�J�*A �����6fg��$H�"D�:�
�'B���N�h�
(N�:t�Ҭd�/�	�&A���2dɓ A��]]]���!L��*J~���M�˅0�H���bE�җ �a��tܰ�t7_|����XK	a,%�����*̮z�/1=?TcWW= �FD�%�����]��2>>>>>>333+��:t�(P�B�
(P�N�:t�ӝ:t�ӧN�N�:t�ӧN�:t�ӡBѣF�ӡBѢt�ӭZ�jիV�Z�jիV�X�bŋ-Z�jիV�N�
�֎8�8�8�8�8�8�~����߿~���-q�2X�c��߿~����߿~��4hѣF�4hѓx<�*��ӧN�:u:t�ӧN�:t�֭Z�IR�P�hЙ��,�t�ӧN�8�ľ+��N%�լ��B�K������UD%Z4NѣF��N�jխ!B�
��'N�jt��*t�-,Z�;D(I�&L�2dЉff�� @��J�*T�T-4N�:v�!Bt����h�
��@�lϏ��j���������jjg��秧ꊊg��i�	BϾ�&��N�n���Cro�nM�(R���!at����$�a�f�aXV�J&�)4 "HTcHHHTTSSB�	S�D�f| $�R�J�$��*LIT(P�B�
(P�B�
�ӧN�:t(P�B�
�4hѣD�ӧN�:v�4h�j�(Z4N�:u�V�Z�jիV�Z�jՋ,X�bŋ,X�b��d�c!�q�q�q�q�~����߿~8�8�~8�8�8�8�߿~����߿~����ѣF�4hѣF�`�h��&L�2dɒի�Z�b-4N�;F�֬dɖ�9ӫ_�X�vKS�ZѢ��#�N$�!�#d�;!�-ht�֍!Z�j���4:��u�Ӵh�
��2B�:թ�!:�D�V�N�	ҢI�:t�ӧN��Ʈ���b�����@�� @�"D�*t�֍!Bt�ӧJ�*$H��D�B��bN�BtI2dɓ&L�2d� ���~�L�7�4�&%�N�� ����CB����K��FF"DA]]]���! �2�8x ����w���C��
K.�s�PP$$$81�  (.buc!"D�$H��J�*T�S�N�:t���ӧN�:v�4hѣD�ӧN�:v�4h�j�(Z4N�:u�V�Z�jի�Z�bŋ,X�bŌ�2X�c!�d�c!�~����߿~����߿~����߿F����߿�ŋ���4h߿~����߿~����ѣF�4hѣF�q�8�P�q�,�����~;�ߎ��&K,d;��q�w�߿~���L�-Z��!�q�q�-Zɒքʝ:TI�(S�d�:թӧN�:իV�Z�jիV�Z�jխ4N�jըP�Bt��"J�:�F�Z	����{15u61(_� $�1*��RZMj����	d�:eD��h�	RbN�:M� ��䔔������`5��t������8Ȉ (P#���
�x�=@��nh�l�˫��Mk�1�rXd�����_��UDl7��3��J��l!����v���`�,�*T�R�J�B�
(P�N�:v�4hѣF�4hѣF�4N�:t�ӧZ�ju�ӧN�:t�ӧN�jի,X�bŋ,X�bŋ,dɓ&L�2dɓ&L�2dɐ����8�;��߿~��4hѣF��8�;��߿~����߿~��4hѣF�4hѣF�4hѿd��얡d����q�q�q�q��%�2��8�;��߿~��&K�Xɐ�8�8��d�kBeP�*$��,Z��t�ӧN�jիV�Z�jիV�Z�j֍'N�j֍!B�B�N�hѣF��N���1'H+�:Ѓ3�U�N�h�\J�ĴZ���Q'P�N�	���7Hh�srk�*+;;;;;;;9IIIIIIIK��� p�C �a  �1�����w;��W��1%������ca�B�����$9�X�x� ��������@�O���O�S������221@@GH����R�J�*U
(P�B�:t��4hѣF�4hѣF�4h�:t�ӧN�:t�ӧN�:t�ӧN�:u�V�X�bŋ,X�bŋ,X��&L�2dɓ&L�2dɓ&C�;��8�8�߿~����ѣF�4c�8�8�߿~����߿~����ѣF�4hѣF�4hѣF:��V2Z����X:7�߿~����߿~���L�,X�w�8�8�߿~����X�jՌ�q�q�X�k&KZ	:�	Q'P�h�jv��N�:ի-Z�jիV�Z�j��S�hѣE�V�NѣF�!BѣF�-N�:ֈI�B�K�3�U��Y��#
p���
�&T��bZ�T���h��$��'Z*t��ӿ~������������(ַ���tJ-���G�n�����\�G~����������qs������ѡB�k'�N�:t�ӨP�B�
-4hѣF�4hѣF�4hѣF�ӧN�:t�ӧN�:t�ӧN�:t�ӭZ�bŋ,X�bŋ,X�bŌ�2dɓ&L�2dɓ&L�2q߿q�q�~����߿F�4hѣq�q�~����߿~����߿F�4hѣF�4hѣF�6KZ4Z�kFOߎ�`�߿~����߿~�����2X�c!ߎ8�8�~����ߎ�būV2q�q�bլ�-hUD%D�B�:ūZ'X�:t�V�X�jիV�Z�jիS�N�F��Z�j��ӧN�:t��4h���P�|:���"_AAO�.��#��JM	Va,gJ���T�V�_�ɴd��;������߿~����߿~�:u��~���;&L��3_Ͼ�䋵�e�U��|\Z���F:֋Y#F�qߣF���֭��X�;E�,Z�j�7�B�
(P�B�
(P�hѣF�4hѣF�4hѣF�4N�:t�ӧN�:t�ӧN�:t�ӧN�jի,X�bŋ,X�bŋ,dɓ&L�2dɓ&L�2dɐ����8�;��߿~��4hѣF��8�;��߿~����߿~��4hѣF�4hѣF�4hѲZ�
u��~�u�F����߿~����߿~ɒŋ�q�q����߿~��&K2d�q�q�2bլ�-h��v�D�B�bŋV�d�:t�V�X�jիV�Z�jիS�NѣF�֭Z�jթӭZ�:t��4B�KE�Z'fBt�0�(_�K��ޭŬ�"�����%Oŝ%��оBA����ɐ�߿~�����~;��߿~�������닝얧X���)D���ī��Y��a�s�q�Dm�ŭ�B��ŨP�Z�:իV�Z�jt�V�Z�i1-4|W �
(P�B�
(P�BѣF�4hѣF�4hѣF�4h�:t�ӧN�:t�ӧN�:t�ӧN�:իV,X�bŋ,X�bŋ,Xɓ&L�2dɓ&L�2dɓ!����q�w�߿~���hѣF�1�q�w�߿~����߿~���hѣF�4hѣF�4hѣj)�;'��X�to߿~����߿~����,X����q�q߿~����߲dɓ&C�8�;&C�Z��%�'N�蒧V�X�:u��N�:ի-Z�jիV�Z�jթӴhѢu�V�Z�j��V�N��F�N�&ёV���Wc:�i3�pb�j��k�=x4PX�l�RZz@�IR�d֎�����X�bՋV,X���L�2d�:v�!B��ŭ
�|WfWH?/%"Ty�$����ֵ��#�0j(�������X[��]�QL������y��꺻3�ɾ>> L�7��gD�:��ӧN�:u
(P�B�
(P�B��F�4hѣF�4h�:t�ӧN�:t�ӧN�:t�ӧN�:u�V�X�bŋ,X�bŋ,X��&L�2dɓ&L�2dɓ&C�;��8�8�߿~����ѣF�4c�8�8�߿~����߿~����ѣF�4hѣF�4hѣF:�(S���!�b�ѿ~����߿~����߲d�b�C�q�q�~����߿~8�;��q�q�-Zɒ։֭NtIS�4Bt�u�ӧN�jŋV�Z�:իV�Z�jխ4N�jթӧN��D�Ӵh��ҭ
�c&��PĔ�֏�n�8�e�-�YU�0֠��ܬ�3Q6}9^�JdʓfHH&L�2WWWWWWWWTTTTTTTTfWWccHTTcT=#"
x ��D�8�5�5���6�����>�DDG*l�i
��j�όjjj��Ϗ����� @H��V� T�S�J�*T�R�P�B�
(P�B�
(Z4hѣF�4hѣF��N�:t�ӧN�:t�ӧN�:t�ӧZ�jŋ,X�bŋ,X�bŋ2dɓ&L�2dɓ&L�2d8�~8�8�����߿~�4hѣF8�8�����߿~����߿~�4hѣF�4hѣF�4o�4B�th�8�����߿~����߿~��%�2��8�;��߿~����d;��8�8�Z��%��Z��'N�:$�4+S�N�jիS�N�:t�֭Z�jt�4h�:t�S�N��F�Ӵh��Q$��9S|"S%P��r���3� �����M�P��J�'��M��$ɟ�����*$1��������*********)�����������ȟDd���!P���'�a�)��kk�T�hd�\�ڒ�2~FJ�#=999/=Tcf|||fff| ���̮�������@�1& `��P�|*T�R�J�B�
(P�B�
(P�hѣF�4hѣF�4N�:t�ӧN�:t�ӧN�:t�ӧN�jի,X�bŋ,X�bŋ,dɓ&L�2dɓ&L�2dɐ����8�;��߿~��4hѣF��8�;��߿~����߿~��4hѣF�4hѣF�4hѿb��Y����7�,d��8�;�L�2d�w�ɒŋY2dɓ&L����u��~�vK�B�u��NtI	�*t�B@��Z'*%
v�N�h��F�� %
(J��?"Z�:�/�ӭ:��E�X�IA�H�@�H�@^�C�b����z�y�K��jd�������|�l0;!Li�>��S�H*u �M�@��2�Ae�&/��FFNX��C���LA�T�])��2�"yJ��ǆGF���

���H������@��NX�ID�������+� ��Ʈ�^�@�31�����*~�	ҢJ�:t�ӧN�:�
(P�Bt��'NѣF�4h�:t�ӧNѣF�4h�:t�ӧN�:t�V�X�bŋ,X�bŋ,Xɓ&L�2dɓ&L�2d8�8�8�8�8�8�����߿~����߿~����߿~����߿~����߿~�4hѣF�4o�d�j�C�u���얭d;���q�dɓ%�2d8�2Z�h�8�:1�����C�8�?Z�`�S�N�	Ro���ɾ)��BU�A$
�:T��(P�:TJ�����es�bQύ��	:���M�U1Q�pB"0@�2!G����D�)Rsgn`]P`UEV2- U55@@8888kRg.>@Er��B�ى��Uē&�FrbL�����A5G�c�G��Ay)y��){@�X;�,�XT519���%�JR_5� ��$�������B�H�������������HWTS|fcfHf ��@�R��D�h�t�Q"D�*T�R�J�*�
(P�Bt�-4hѣF�4h�:t�ӧNѣF�4h�:t�ӧN�:t�V�X�bŋ,X�bŋ,Xɓ&L�2dɓ&L�2d8�8�8�8�8�8�����߿~����߿~����߿~����߿~����߿~�4hѣF�4c��b�C��q�,d8�,Z�c&C�8�2d�jիV�X;&K-Z��&L�2d���?F;%�,X�b�IЭX��t'N�̨~��̐zz�L�C���	�ff| A��������yyx8Q�y����d�Dj��CAF@���ǋ��,
0R��������ܪ��j�R������������|�|\�ld��z���$an�v��$
�����HHS/H/ST/#9#"})���������LQW�Ji}��°ċ��QkL4<.6636l�[%� 0�p!a��Z��(�)�y�1���A��bɳ:L�ҩS�*$�2dĕ*T�R�J�:t�ӧN�:t�ӨP�hѣF�4hѣF�4hѣF�4N�:t�ӧN�:u�V,X�bŋ,X�bŋ,dɓ&L�2dɓ&L�2q�q�q�q�q�q�~����߿~����߿~����߿~����߿~����߿F�4hѣF�6L�2d8�8�,X�jթӭZ�q�2d�bթ�4h�:�K-Z�;D�ӧN�:q�-Z�vKV�NѢt�S�&���%D�*T�����������Y���OO���LR@��H�B�`�@���a���FNK����O�B�AC�@^a�QbѦ�K`9��������������������������p�j���\pphd��Z�)kw�+� �}"�Aܤ�ii	j���6d���53�s�Ps�1P7ӥ�p^E�F�n� �"4BP}�ĕ�|Iv�ǈ"�������l;�����jg�li!o�eCc�$�Ć2��d�ٙ�ʡ&A����2dɓ&L�2eJ�*T�R�N�:t�ӨP�B�
-4hѣF�4hѣF�ӧN�:t�ӧN�jŋ,X�bŋ,X�bŌ�2dɓ&L�2dɓ&C�8�8�8�8�8�8�߿~����߿~����߿~����߿~����߿~����ѣF�4hѣF�jŋ2dɓ%��hѣD��4h�bիS�h�	ӧN�h�:v��:$H�"D��:�V'B��ҥN�BU���6evg�ɳ$�����������|T=?S?%##99#%}���>�EDA�@�Ȃ��AT��@B�AB�A�B��C�F]�/Ѳ�x�[#N�iJ�#�۫��S��Z�R��ꂂ***�zZ�*��
Z��z��sQE��l��6���@F'�Ag !�$Jj�G"��,d�����\ŲnD$z!�aa#x5�p��4�@��AQv����Dܥ/�ȃJ'�����$<��z~Fb�z~�Ʀ�ƐƮ�bz�U ��f3�����τ| �A��dɓ&L�3�N�*$�S�P�B�
�4hѣF�4hѣD�ӧN�:t�ӧZ�bŋ,X�bŋ,X�b�L�2dɓ&L�2dɓ!�q�q�q�q�q�w�߿~����߿~����߿~����߿~����߿~���hѣF�4hѣ:�:ŋ,XɒŉН*uF�N�Z���D�:TH�"J�h�	ҥD�||||||||BtIT-�*$�31"_�����ٕ���NLLLLLLLLT���NLOLNK�K�H��_G'$��b��c$@o��S�<��,<<TD<��z�������Fð�i��l��=��9���:�&��000//.����7�����*� %����&59����*�����6�^cnǙkr�hQ�xs����
	2,x��;U���,3�6pD%�D��hdx֘|����r��I�_�y�7���E�l��y���	@�A�Lj�F)�o�ɝ�MiT�llillτ @�
�$H�$ΡB�
(P�B�
(Z4hѣF��N�:t�ӧN�jՋ,X�bŋ,X�bŋ2dɓ&L�2dɓ&L�q�q�q�q�q�q߿~����߿~����߿~����߿~����߿~����ѣF�4hѣF�IV�V,Z�b�L�4:$�S�*M	ҢH>+��L�bD�*TI2��������� @IQ$	�1�$1�WS=HcS?SHTTSS??=1111==/9/??9%/1//999##}��Ȉ�C$�d�$@b�O��0�0pp��P�xk�0$P9��p� =#N�Ô��I�III�՝����������yuyy�AUA@�U�-Y%U5Y�@� ����Y$����Yu$ѭ���Z��|R0�dހf!J)Wj�A(f��C��!p+��Тh��ddd�ꊔ/�nR��Xg����,05�\��($����� ��A�DU����
�+�***$+�>33333333>>>>>>>>*$�2:t�ӧN�B�
(P�hѣF�'N�:t�ӧN�:ի,X�bŋ,X�bŋ2dɓ&L�2dɓ&L�8�8�8�8�8�8�~����߿~����߿~����߿~����߿~����ߣF�4hѣF�(V�X��Ō�,hT�'P�:$�Q$���� ��@��"I� �����������M��2�����������OOO��LLLOOLNIOOH�G&%䤤���!P���<e�J*r�9l<����FAȀB��A@�b���0��g`p`б� �x���CCH���6˰���������թ�I큹5YAyՁ��@�-uuyu���5y%�Y�%���- �YAT�U-��k5a_q���cu�Av��!}��FėC��XW��0�%X��Тh��Iv��$@��v�����	|�7�gj�����F�"¨����biKqH@�q�(Y
jjjj��l���������������J�@�N�:t�ӧN�:t��-4hѣF�ӧN�:t�ӧN�jŋ,X�bŋ,X�bŌ�,dɓ&L�2dɓ&C�8�8�8�8�8�8�߿~����߿~����߿~����߿~����߿~����ѣF�4hѣF�@I�'D�:�jũʓ �����������������@�dɓ&@����vg�����������li							lli
�jg���������	
�g�&&&&%��$ddDB�DO�RR7�蔍�*JzF��-""w��<ޢ�.�s���w;��7s�X$81�� x�����Õ��l���)"9����������&���00//(((.���/(/00.���(7��.�������59�� ��_Ͼ7+�Ð����k�	Jpr2B��,2�7F�Ap	*'��	m�A��K�x�P����������A�;
8/(1�a�Ǝ#g%�t(�\�Y�Ic�-�y^&%�����s�00��604)�o�Ĝ��fN�u�řb�3$�����&$IS�Z4hѣF�'N�:t�ӧN�:իV�N�jՋ,X�bŋV�d�bŌ�ɓ&L�2dɓ&L�2q�q�q�q�q�q�q�q�~����߿~����߿d�q߿~����߿~�q���IS�I�u�խ� @����g����������&L���ٟ ����̮��Ɛ���������Ɛ�����������~���~zb^^bb^^^rrFD*D�%%%%#}����
��>�a�$DB�b!�N���!qGs���y��o7���(�w=E�C���� �а�i��l9\�W+e�ZR������������������������������ܺ��R��Ԥ������z)<��nW��&��>ᐡ(��ܛ�{<�ȟ|oaXf��J*&�&��

�
��O��}ӴG ��yJ	Q��!J�n��\���yD%K��:�Q[�XP����a�5����P	����T�] �QQ	�j�l��:T���zu��Z4h�	ӧN�hѣF�'N�:t�ӧN�:իV�N�jՋ,X�bŋ�X�bŋ2dɓ&L�2dɓ&L�8�8�8�8�8�8�8�8�~����߿~����߲d8�߿~����߿~8���@H�d�>*ѣC�D�&L� L�2�����������������������������O��LK��NLK���NNH�D���ddg'$de�&'$��'�b����Ac / сq�qqqAG��PPPPQ�(((.(�w=^��!!��� ����,v;W+����I���������՝�������5�����՝�y�Hhi��x�)(8�n�JP�A�^R�[�R��ٵ)rO�L�[�
&�&H
���j�ɪǍͬg]�E�.���Շp����<��TB}�ėؠ�__e��QL(���`��2�J�4�����$����e��y���31�	1X���L�5�I��X�ucF�P�:T�F�4hѣF�4hѢt�ӭZ�bt�V�Z�bŋ,X�c&L�2dɓ&L�2dɓ&L�2dɐ�8�8�8�8�8�8�8�8�8�8�8�;&C�����߿~����8�Ϗ� A]��S�N�*TH�dɓ|||||||||| @�2d�������ٟ����������������������K�LLK��NH��K���NNNH���NK���K��O��K�H�\/W�x8�Ph����y�

��������

����
<�oW���HHpp``c���z<^�B��c���r�[%�*JJJJJH���ooonnh���n�-��!k`�t�t�I���y�7F��_��_dP�5R�l	i�c732��!ML�[ۗ��JQP�ae,%�M�(_|Av�"D���+��!J��+�%*Q3(6���J�bH�|ltR�W洫��K-I��I�q�0������4��Y���:L��%J�:�
(P�BѣF�4h�:t�V�Z�:իV�Z�bŋ,Xɓ&L�2dɓ&L�2dɓ&L�2d8�8�8�8�8�8�8�8�8�8�8�8�ɐ�~����߿~���;�����d�ٟ	�*t�R�D�L� @���	� ��̮����Ʈ������A��񙙙]]]]]����]���!QQMQL������^^^^rrrrbbbb^^^r^^^^bbzzzb^z�~brzJ~D,�} �
;��1G���(..000000.......00...�y����s���	 x�^��CN���ca��l�JJJJT��������."�ñ��s2v�J�a҅�܉�]�܈)I�a"�#��g54Qmqk>I85VKI5E^Mj{Rr�[.W)k�9KRf���toF���Qt
$��T�QJ���J+�C�a����E*``�3(>�.%�n��@�P}����$�*|�0�`��n�P�����̨^��@�R�J�*TH�(P�B�
-!B�
)ӧN�jŉӭZ�jի,X�bŋ,X�bŋ,X�bŌ�2dɓ&C�8�8�8�8�8�8�8�8�2dɓ&L�2dɓ!�2w�߿~����߿q�&A��������T�R�D�&L� @���	� ������Ɛ��������@����332����B������y�+��������������ļ�����������������^�t��

<���o1AAqA������qqqqqqqq����AAAAAAAAG����z�8\.���X�x������e�ZZZRRRRRRZZZ�r��!��V�o7.��,"�J�v�	�r�7IT��ਗ਼�M���	���²*�꩑��k:!k���j��j�Jw�l���_}��
Q�Ǝ�7�UŴ��͵E���E�̸�����q3t8�
$��E�`�tZ���j���:\�j�#����JR����b��bP�:t��d�B�
(Z4hѣF��N�jՋ�Z�jիV�X�jŋ,X�bŋ,X�bŋ2dɓ&L�q�q�q�q�q�q�q�q�2dɓ&L�2dɓ&L�2w�߿~����߿q�L���2�D�&@�1"D�L�2 @� @�uv664����5vg�fer>>>33+��������$**)������������������������������������������������
����<��������������� ����� ����n�p��Hp`c���p�<^�B����c���l6�V�a��v;%�W�a5 �}�7K�������7�]������q��Sآ�Ģp|��h�PrXW l�t�+&6��%R�GyS���"o��K���(�(���5������������5����������e�͵�D����s1��lÜ �!���@{��R򺫜��+�$1�T�ӧN�:t�(P�B�
t�ӭZ�bt�V�X�jիV�X�jՋ,X�bŋ,X�bŋ,X�`�8�8�8�8�8�8�8�;&L�2dɓ&L�2dɓ&C�����߿~����8�D�| L�ӥD� @��"I� @�dɓ&L�7�� A]���!!!Q!�]��\��������lllllj��jg秦&&'���������jj������jjg�����jj�jjg�'$d@�!���{��,(0�z���
<�b������������ C�� @A���C�₏7����		p�<^/G����z=�G�p`c�ʬ!7"��f�JXw��_���*�T �y����K	9F�6���7��
�_f�rD$���isaE*�0t%TU�_��'Z���D(�n��E����٬�1���й����D��Dʹ����D���D�|�J�Wė�[��R��$lQ6gUT^0�6���L1�r"*^�@�B�J�*t��(P�B�
�ӧZ�b��֭Z�bիV�Z�būV�Z�jիV�Z�jՋ,X�b��q�q�q�q�q�q�q�vL�2dɓ&L�2dɓ&L����߿~�����qΝ*T��"J�*T�R�D�$H�"D�$�2ٟ|fWcccccccc||||||||&@����f666666664�EE3��Ԅ���EEE55D�664���u3�EE64���3�����P��� �x��@��������������y���1q���qGp����t��������!�Gs���w;��稰s� ��4� x� 8^�G�cQ�%�7&�o0�Նvݷ��$I
P���W�B�/ĸ.ՇLW�6�+1"��\]%Bc��"���k�Ke���Ɯ��'%~��n���JL��؍O�Z�������[[TTTTL��\\L�AEо(�]	R��K���kLJ��9�  7��1�� �����S�f*UM�E����jՏю��&KZ	���V-h�jŋ2dɒũӭX����;&C�8�8�8�8�8�8�2dɓ&K,X�bŌ�;��ߣ~;%��8�t�ҥD�T�R�J�*$H�"D�$H�$ɐ ���@��2� @�2>>>31�����������*)�������$**$$$$**)���+������������A��].��'s�\4\Q��w����
;��C�@B�₂��Q���{� ]��t��<���s�� �,z�� <^/g����,4p|ܛ��%�A����rXg"_��>�6l�r���s� '�h�ؐ��Z��.���d%U'���UV�q���hIw��K}�7EUc�%c��c������cCB���ƶ�����337C���`!(������I#c��UU�爰�#�s�T4�����bU��NЙ��Z�����X�qֲF��$��Z�jՋ2dɓ%�S�Z������&C�8�8�8�8�8�8�2dɓ&KV�Z�jլ�;��ߣ~;%��8�t�ҥJ�T�R�J�*T�R�J�*$H�$ɐ ���@��32��������ɓ&L�2>>>31��������1�����$33+��������)�������1��>>��������<��W����x<��  ������p�k���y���W����y�8C���q��@C�\Q��w<�CCC@����]����, � z�<@�������}�|l�8	I$���&@�v���K�a��j��4��h����J��`�`1*fd��0��QJ������X��BV+>��@k�7h/���R����
����K
	�񱱡�qqrbbc[kkj��������������Y%*Q<V<^.t/���&�	�Fk����e��s s-v<�Y����0�w�*�I�:�N��E���B�jq(Q�*�:u�V�Z�bŌ�2d�bիV�d���ɓ!�q�q�q�q�q�vL�2dɓ%�V�Z�j�L����ѿ��L�q�:t�ҥJ�:t�ӧN�*T�R�J�$H�d�f| @��ffffffffb	�&L�2d|||fWWWWWWWWfffWWWWf||||ffWWWcTSSTcW*�ƨ^~̮~��D�x�]"�7���k� \`Y�X,�y��;�@B� B��������\P\``PQ�,�z���;����!�qqq��qGs�]�,� p��:@��Cd��a��퍌��%(����7\]�����ޫ_�H�RU�R#���D){V5PEKo`D)ujgr����KT�MX��V7��� a��Kat�$�HZחPRUU�X����X�PO�������������[[TTTTJ.���2�A�9�*|��l�Im.<k6<3.6I.0bV3LVUV2t%���͑�0�0t��[��- U��,��:U
r�S�h�:t�V,Xɓ&L�,Z�c&C�8�,X8�8�8�8�8�8�ɓ&L�2d�jիV�Zɐ�~��7�Xɐ�8�P�:t�R�N�:t�ӥJ�*T�R�D�L���	� ����������@�2dɓ&L������������Ϗ���Ϗ��|||ffHHHcWW||c1Tc=?c??1-mv�Ǎ��N�e.V�Hp@����t�
������x��X$\\5�00�y�<ޯQag���\P\`\`````44Q��y����瘸�!�.��Pr\���(\$�\�����y!��n#r�-g+҈��,c~ֿ�CW�CT�'���#ÅdUUwT��֥��cT�f:�:��]�����&� ޔ��ȸ���
J*��ƨLLLLH('�����Ɔ����ɉ�mmmj%D�Fה�Y*Pkkk6kkm463Q.L2..6Q34><6Q46$����R�/G6 ��Ո-!�"J��:���ZZ���֡X�jՋ2dɓ&K,Xɐ�d�bŃ�8�8�8�8�8�8�8�8�,X�bŌ�;��ߣ~;%��8��
'N�*t�ӧN�:t�ӧN�:$H�$ɐ �@�2d�>>>>>>>>>&L�2dɓ @����3������������ A�񙙙Q!]]���]P�\��C�%�1�aA�+��.��F�+�fÛ�9�,�x��������q��сg��i��y�^��OG����p�<�b��@N�����w�;�@��K�4Q��x6�"�l�t:K��	K���k�� q��Kʁ%W��Q_ȅQ�����h�MR��[����P
^�Ԕ��ԗ�UUR��ՍZ��"?�*�!y^��&��G"\�����A�����ފ�ޖ����pppdd�����xx||||lhhh\\\\��k3.A0Lq(��&� �5��$����&5����(�*�����:���[*LE��If�Ǫc���BTH�֡X;%�,dɓ&L�,Xɓ!�2d�bţ�8�8�8�8�8�8�8�8�2dɓ&L�;��ߣ~;%��8�Ѣ(N�:�
(P�Bt�ӧN�:$H�$ɐ �@��$�> @� @� @����3��������33����������ٙ��H�IB��S��R��%�p�a�rDB�\�IJ����   5/.�� 6���P��&��(� K���x�=MRF����J^��+`�1�00�w��CEޠ��ǅėm��6�O�M��D@W��iE�M�7"��G^��ԥ|�7�̓K�Q���7��$�$��6���� + *����&!Zh�Xl�F�$�K���݋�y,�Cv9��dp�������ޖ�jjj��ppp���Ă��x|||llhhh�`hf��\�fhl\h\�xhĒ�x|��l\\�j�hl�d�h����AVQ>@.256I>mL4<P^$��*�g��.�m��61eF�	��hujŋ2d�vL�,d�vL�,X�j��q�q�q�q�q�q�q�w�߿~���L����ѿ��L�q�h�
'N�B�
(P�:t�ӧN�$H�d�| LH�d @�	� A��� A]�����>>>333+�1������[�J%�`1���*�"�U��o+�ฺ
(5�aXaoJA�1�(��1��6a�q�����@l6}��%�G�N�I!t8)Dܒ �3B�A�{9K`hh��� p� <S]	R�@��J�\]-g��	/����ݣr���p�Hh���%E�Men{U0=Fx�L>m�	"}�mbJ�nK�6t*�%�$�2:`��ip0�d�aA��f�$�k��� E͆�V����V��eecSST����&$�����cccG�GE��V&�CF�cc�B����c�&�Aq��rbI��q�Y���a��
jJZ	q���d�;0P"
���� U���*�2�u��d�q�2X����2d�būGq�q�q�q�q�q�q�q߿~�4h�2w�߿~8�2d8�;F�4hѢ(P�:t��J�*T��"D�$I2d||||||||||| @�� L��d����	�M����]�QM�P�,)��ڕ_/�.��Zc�*��(%J+�H�l�&8��۶�\��R7���������k�.K��+
��)I�o��"ð���aR��o�D�7��}��.5Ł��||�f��f�%��h��֢\d��då�	��H#q�n2�`�U�d$��I$�/�{򡉪'�++3��/"��:��.�=�5=Md�ج�⊓'�WRJ����� ����W�}��&�w6����5U�TTTT��UcS��$�&&$����cccCccccccccCB�Cc�$�����&&&&&&&&$��������Se�U2'�����:�	=B�r�0%FC�-�;D(V�I�X�
�Z�֣F$yU�Ӳ�N�c!߿~;&C�;%���d�4o߲Z���KY2dɓF�4hѣF�P�:t�ӥJ�*T��"D�$I2d� ��@� @�>>>>> @��$�2���	�|Nu�P�!��3�P�u%�*���ff����\\`Q33(��L
)T���̒!���a��PPW�J`c�༮�1�y^W�r\��a���k�0�KÃA�3
°�+�0��h5)p\���J������ �llP��(�Ά��D����9���Ay!�_v�08!�c[f5pJ$���*��#��hx\|f�/���[���&�FGK������D�9RΡk/���k��@��q���q>�nX�/k�o$�Wb���ꂂ�+{zZ����JJJK
	�������������������K
K���������񢫰P1�,��6Hv7)�x1��6�>>-Z�I�l��:�u��P�XUj�i�Y#�X���Z4Y�d�q�d�jŃ��&C�F����q�8�ѣF�4hѣF�P�B�	ӧJ�*$H�"D�$I2d� @� @�ɓ&L�2dɓ&@��"I� T��1"I���>3+��=�J&����ɉ�mmi�Ɔn-��&m�m�&&fͥ�@�I$�Fͩ�+ȍiRIA�}�������c��+��.��8��,;ø�༯+��+��<�� �p���|�t/�ˍˏW��\i7v_��K��C'ٲ002���o��)�E*�m((F0�&ʌ��&��/50O���X�T�O�ZՓW�SW�U$N�(�]�K��7ѐq�j�}�P��K�<���%8.������������V��UcT��##$���&$�����������Ã&$��T$�&&$�&&&&&&&#########���������$�V�T��aA�Ub1!�n���5�����c���HC2�1լ����Ghtqӭ=&���h�2d�q�u�V���Y24h�юɓ!ߎ8�hѣF�4hѢ(P�Bt�ҥJ�$H�"D�$I2dɓ&L�2d�| @�2dĉ$H�"D�M�]!P�31�*����ȦMff�G���ƅ�ɉ(&�meɍ�i�ɍ�-eǅ�n�A����Pm<2ME(/����D��0_%R�����>�a��B!�۶�n����B6>ϰ�lI0qt6��S[MO����EWn�	�Ky~����SpaT�Lc���/�"�TJ)R�Tl�8�Ĉ˙�#�kp\aD��\��%)J^RJTl��	����YE\���ɨPb}�ѧSa؅E��qJJ�/��f����+��Q]Yڛ�XWT[��U�MP�RRX������������U���PPRՐRX�RRRRRRRRN�QP���L�[-�e`�1Q��yc��A
�����6Iġd� �x��Z�E�.u���"e_��-�7��2���2~�j�ߎ�c!ߣF����X�bփ�8�4hѣF�4h�
�P�:t�R�J�*T�R�J�*$H�bD�$H�$ɓ&$H�"D�$H�$&L�332����H1���ɉ,H(,LG��LH'��Ɔ��G����ƅƆ��mf��Gɍ�mm�+��&tS7AE�``�����tJ+�$�P(
����g��}�gؠP(	$�JU*�t/�
&�$�ĸ�1�����$�Y��%�a{���y-�v���;g����GC���oɯ���1v��QUk�7R������aA���}��5�(<�H����(�㐥Ȉ)IE!L����S�h�K�����7.@r6_���!���sp��))"9���77&�/.�"�����++��� $����������$�11%���$���                +*�$� �1 ���!��e���B"��@b��n�WK2!g�C��d%�p�})���6Y��=1"t�����Z�c���~��RkS�h�c!�,toߎ��7쟲*8�ѣF�4h�
'N�*�	ӧJ�*T�R�J�*t�ҥJ�T�R�J�*$H�"D�L�2dɓ&Ʈ�$�Q"D�T�6e5r7{e�и� ��ɉ�%%%����X�%����ظ��������1��Y||f����ڢf�ff�`�t:
%��|�J�W���D��t:
%C�������Ŵ̢`��x�|l�d���ꚠ�7NA_���o! ��M�H�%�!Cl��;d�A��q-���B��|l�F�DU�~$O���Z�LX��Q�����
%�v���$���Y��J�e�����k��!aa CrH��)@�۴G#Ez��[%*Nol���ɬ˪���ij����Ʀ�����FI)*�ƧFGFH'�Ij�'�H'�F�g�.`
��).���b�$G�@�3����5Y �t���1�,���!�˚��x���f(V�NML,��\J�V-Xɐ�d�6L��Nɓ&M4hѣF�N�*T��(P�:t�R�J�*T�R�P�:t�R�J�*T�R�D�$H�$ @�
��ό��
�
�	����.��#�TT�$��Uc��SSTD���###$��#V�$&#�c���dDCc���D�����ƶ�3375����ֶ���ִ�����eU��֢���)J,"¹�I���k�r 5HP);'���Z�܍�VwAs��fڢf��.6}�OϛNS��I+���5�QA6625MsjoK`uV.X�Iy�����e�ѡk5g ;�J\�q��n]��D��)@ q8.���Ô�I��՝��5�yuu���--UUUYX����-Y ����� ���� ��������� ���������$�ىY �� �% �$�%�Y��٬��U���8<Q1�� Π\x��j�\|��� {^@6<v�6^�P�|9x3�����	:�:Ռ�,Zub���,X�cF�4hѡR�J�L�'N�*T�ӧN�:t�(N�:T�R�J�*T��"D�L� @�2ʅ�C!�HS�a�Ԭ�������jp����p��jj���ފ�Zނp�d�pjj�d�p��jp��dd�xx�Z�QLK.bI22I<4L<<>644..LLLkkmmmQQQmkL....446666>A>4AVU2<5EE]u))V}����x����q9��Ix���, �q0<4bx!du����Q3LyRGd�1$
IA1Y�E�a��F��K�64I66@ogR{MPU2b8;��Kqb��F��ږ�|��jz�M�n7h�����(M��(��F�44�l��9����7&�/.�(("����������++�����������   �         �$�+$�1$���$� 0  �&&�%�;�NNR�RL�PQ\L�QZ̜.T"H)��U[SAO��َ�N�b��Hf%9:��իV�hѣF�!B��ӥJ�:t�ӧN�:t�ӧN�B��ӥJ�B��ӧJ���@�2gD�+�>>+��3�F��[������������������������U�T�WK[��������R���[���L�P�JF�O��MMP��PO�������������L�P�����P�]MMUZ��F����_��xމy6 D�n���� /P�A��(�6� (�V�:�`|h���QK1B"@t�K$����`c�_po$�Xd�|�!rD#d(�j#R��#��Gr4j�DK�������Y�7�f�v�o9~��_��t�sy����׉j[�͹�՝y-AAA����---UUUUY ��YT��������������������������-E�����������%%%%%%%%%%%T����ɼ�%YUYU%%%%%%%%��%���4(���t���� ��N~"�ѣE�U��W�GZ@�$�4hѣF��Bt�ҥN�:t�ӧN�:t�ӧP�Bt�ҥP�:t�ӥD�&$���3�F5uB0�'��`��-uuuuuuuu�A�y�5���������޺������ޠ�j������R�dj�����j�dd���������Ă��xxxx|||xx�����xxĀ��|���������}Ӑ\��Bo@_�@�Jȴ$8�� ���5�d��Ef�U���R���h¨`���F��)m��)%�7���(��.K��kj1�\�ap0l��IF��%X��DFȂY�I���T�ޗ�yW��7"
�.@7����4�^^ju{un`]^PPPPEEooKKKKUUUV@@@@@@@@UV@22@VU8888888822222222IIIIIIII2bPn8<2AAAAAAAAA<<<AAAbbAAAbbIIIIIIIIIIIA6>I2bI@A22bAbIb88888888IIIIIIIIAbA2I<R"�M8bbLbb=t�QP�N��0� Qx��C���4hѣF��Bt�ҨP�B�
'N�:t�ӨP�:t�R�N�:t�R�I�> ��̐zF2�l&��9����////////////////777777777&�75&��X��TY���W��[�\�ڗ[�U��[���U�MP���RRRL���R�MR��ے�]��DE�_�ݦ��Ar �/��v�4r.�;���D��1ш�,�u�e泃7A�i�E�Hޔu������w�D_�~���_�nv��_����Ⱦ��HM�	v�I"�/$aީ��rw�����T�#Tcc�g�rc�&���t�.bv�I�0͑F�qJ#�s�򂂂**+{zZ�����������������������������������������J�Qᡑ������������



JJJJJJJJJKZ�Y���
�J
I�JJJJJJJJK����K�����0���{M2>,Sc=83A30v$-*��!ͣF�4hѣD(P�:u
(P�B��ӧN�:u	ӧJ�*$�ҥD�%	4�5Er�DEވ�����ɩ����������������������MMM�MMMN���-MMM���MML�LȊOl��ȫ΢�V�Զ�����TTV�����������UUeecSUeeUUUT�e�w6u����*U�܀n1�9�7F� h;K�<����A �T�D�'��

�'J��ў�1��L��#82()ƚ�\K�e�iE*��P_8 ѱ$B!(�5����1Y�Ú#&"�sqoUA���� �5�=Kl��XV��_���E�JE���p����507���������+++��         + $�� +$��������11111118�9� 1 ��� ��111$��������6��1 ����&$��$�1111111111111111$�6K�i��))'���hɇ�����񱡒��(8�[��1�F�4hѣF��:u
(P�B��ӧN�:t�ӥJ�$H�"I� @Ifg�d���'��rksSs;;SSSۛSSSS;;;;������������;;SSS;S;�"#���;S;���;�Rk:�#SSs;�R��`c���jjjk����������ꂂ�*+z***����z*���S��hc���7� ���<��7N@_�l�+�����C
�!i�/5�%�� ���.��X��l�p`H��X%�:�A�4�7�d�D�lj�S� Ubv�V-Z���t��*�`�%�Q�EAUb82820-:A���o�7XK��_��B!������Ԛ������ޖ������jjj���pp��������jpd��dpj�������Ă�������xxxxxxxxh�|�Ίxhxxxxxxxx||||xx��xxx������������ĂllĒxxdx�醦�lH(((((((,LLLLLLLG��LI��!I�����H�%�lG�,N�6��cDķU�U%�V��F�4hѣF�!B�F�4hѡӧN�:t�ӥJ�$I2d� ����$K��;�ʤ�������������������������������������������R���������������Z���������n^nnu)jjjjjjnnnnnnnnnnMMM```^^^^^^``MMRsgjuRl�[�Q�@+�<�H$v���ޒ�(]�H'h�j�AG=)0t"��(+%���*�0�b��`��('笯���#x;�A^�E�B��H�xX[����C�Q�..֓%"gIB��Y��jK9��A��È�>���9��O�Û��nAIojjE@5KVVVV55@@@@@8822222222222@8IAAI8@AAAAAAAA<<<<<<<<>>>>>>>>kbAAooA.>>>>>>>>66>>><<<><<<AAAbbbbbbbbb@bb2I>6Ab8�h&�((((((((((((((('	&�ǉ��)&�&ͦ�&��(((&�ɇ�ͩ�'�-��*Ǝ-f�&�&4hѣF�4h�
-4hѣF�N�:t�ӥJ�*$I2d ����Ɛ~^�suguuun`ugu{s{ujssssssssDDDDDDDDDssDDDDDs)DuDl�9��������":���
ST����CEƚ�]T�JZ��ڙ�ښ�����ښ��������SSSSS[����WW�ƞ��N&����7�t��7sv/��[�\� N@v������6F����TU�V��V���Ȧ���SS�hY#F~��	��8���W�v���e��A_��;Aȝ��ݩ!}��o�-�j�댆_�~��Ko�WV484>46.QgB�~��pj��ܖ�d�޺��xx�nU88@@@@@88822888222IIIIIIIIII82bAAb28<<<<<<<<>>>>>>>><<<<<<<<48>L226b>>>>>>>>666>><<<>><<<AAAAAAAAAAA8bAIb64<<66b@@@5AAAAAAAAAAAAAAAAA8<4b>>U8L6I4L<6mL.<b.mkL@5.kbbkL66>>L4V.2ALhѣF�4hѣF�P�hѣF�4:t�ӧN�*$H�"I� A���]\�d` ��Aթ������쥲�)DssssssssDDDDDDDR))R)))))Rl����9Z��J\��%��▦�7���e͹�I��DgggguuuguuuuuguggggjjjnnMnnnjjjg{guRs8rXE���.D�A��k�ӑ���;	,%|F�\�jjܬ޺������j�j�x2�J�PrR��-���f)�F������ON��<�0�<����F�FM�<�_��|@݄�<����O%�ݎ��@^M��u��ӎ�e�.�%]1%0�0��Ij%r��l���aQ,�:�єU�USÃ��#$�����#$����&&&&&&&#�&#��##�������������������������#$ƶ"��c��������ccc����������#��$cDe��d#C##B�f��#d#C#�C�#C�#&$����C�D���V$�&���իV�NѣE�S�NѣF�4h�
�!Bt�Ҥ�>3> �Ʀ��Ɛ~"0�DsDsuDDDDDDDDRRRRRRRRRRRRRRRR))))))))-----)))l�JT���J]KK���*NjH���+;�`i���0�μ�XX�Έ�������������戈�������������Ԉ��g--p^H NA7`��҅�\��v���^$�!�7��߬f"KkKK`n``MM`]PE^K@Ij>
~��B�.���'h�bw���7��6nуyO!^N��v�v�7�ox�k����_w�@�y0o ��Ar�L!�M�OkJ�F��Up�+"f�)�ͬ1�D��J8�P��z�uQ�;2{%�έ<6K8<2IIIIbbAAbbbbbbbbAAAAAAAA2E<AA6V><<<<<<<<>>>><<<A@L.<kk<>AAAAAAAAA<>>>><A8L6I6>2I42b4>Ab2IIIIIIIIAAbbbIIIIIIIIIIIIIIbbbAAAAAAAAAAbbbbbbbbbbbbbbbbIIIIIIII<<<<<<<<bAAA<<<>bbbbZ�jt�4Z�:v�4hѣF�P�:t�ӥJ�cW| A�]!����L�=��l9��6J^�
JJJJJJJJJJJJJJJKKKKKKKK[-��e�ZZZ�l������Q�JQ\�#NW(�Ѳ��� l�C��)K� ��ʚ�����椈��������������������������R�,$�[�49�RZ�������w��d?f"KLKK`n``MM`]PEPU8bn4x2d:	�@}��'��H1%cx�����<�>！/�y97��o1�~����%���@^ND�:�k�A/�$�CtYMEB�	�px)¦��C��0��}��G:xE�25ƇV�Sf�2�hl�lh����Ă����������Ă���������x�xl�xxxxxxxxx||||xx��ph�ph\�Ă�������Ăx||x��dh�jx|d�xd�|x��d����������Ē�dddddddddddddd������������Ē��������������Ē������������������Ă��x��Ē�j���4h�:t�!BѣD(N�*$IQ"I�&������ƐƨbJ2�p���59�[�e%%%%%%%%��������W+e��l�[-�+���r�\�W+���-l�\��+���r�[�h��c��X�x���h�����pqhs�� XZΤRZZ��RR��������RR��������������Έ�Vzd=q��ʲB�WZ��qV��������V��S$�z�M,1y��8L)X^�Ò"��%<�o)��o5���u����������)����y����7��I� � ��n�����zP}% 
2�B ���R55�v�J��Q(_f6K;|?WQߴf:�����0���%����T��������������$���$���������%��$��YA$�%$����%$�$��������$����������������������$�������������������������������� ���%%%����%%jթӴh�:t�!B�
�J�L�||||WcHHcHS}��)")6[�ײ���������e��l�[-��a��l6��ca��l6�c���l6�+��444�v<^�W+�i��l�@DT�Z��/0 ��f�icд���-r�*JM����������Ғ��%%"�%%$G777TF�k���$��z5�d�ÏQ��$k����W�W���T��NO�\@�#?2-:�p^Pk�)1.&�oE������7�� ���B���7�o0�i��{�'�Ѯч�ټ�yo'��C ��������M0�7Ai@^�ؔ]{��/X�Ģ!(� �A��l�r�j���QF��BU����֒�|x�d||xxxxx�������������������|��|����������x�������xl���|dp��������pd����dpdĊ܀xdd��d��p��pppppppppp��jjjjjjjjjjjjjjjj��pp��������������������������������jjjjjjjjj���pppddddd�j���4hѣF�P�:t�Q$ɓ&��������@�f52�Q{����RR�l9\���d���r�\�W+���l6�V�`i��v;������CCN�c���v;V�����,z<F��Z����d�����l <cE�����jOF�e�4�sDr�K[-��e��---)))RR))RRRDDsr���)3'~�bt�H~F���!Z��Q�SULKUEPEPPPEoUV2II6K(��#9y��)E�$�n��6��j����oB�����$�3���yf��B��<�/�y<}�y
o0��W�'��&��_���$��F�\�ˋ�7�@��Wt�5�$��qzƇJ�h�(]+Yc"O~�<�ld�x��ll||xx������������������Ē�x�Ă����������Ē��dddpxh��dxpd��������j�pppp�j���ܪdjp�l���j�djjjjjjjjj����������������������j��������������������������������jjjjjjjj�����jjj�����j���4hѣD(P�:TH�d A��񙙙]!]�L�(\ ��RZZRR�-))-r����a��l6��CN�`���`�aaaaaaa`�aa`ӱ�444444�l<@/A�˅�4�P5r�@��K��`K���x�)=@T�����c����ZZ�l�[-��iiiIJ���IJ��"""""*�k�sx��H߲G~��1�9r��������V�ST�T����Ud�$��ed��늇�4�|(>�Kz�����[&��o�n��.I"�_xn��P9�nI��� ;@���ȼ��}��7��%T�&��~8���ԍ%Q]� �b��,��
,"�+�B*V�h���q�	�i����JKJJJJJJJI�*	��J��������������������������������z�y�Z���zZ�ZZZZZZZZ��Z[{{{{{{{{{{{{{{{zZZ��{{{{{{{zZZZZZZZZZZZZZZZZ����������������{{zZZZ������իS�hѣF�P�:t�> @����3332B��xhqcd���l6K[.W+e��,,,,,z=�G����,,,,,,,,l6��c���-r�<\ A��Ű4�jR(�nl�
��;%�����Dv)�9[��%�%%%����%%*JJH��JJH��nnk�nR��*k�fȩR�_�d��h�)B=:2�`'
&������ƨI()&FƤ���d�(���D�O��x�㐈	���I nIȒ��_y���^E���@W��r��� NA�B�.�ژ��ù/�D���%�v��vڌV�&$��A(�c�vd��O��������X�L����������RPUMMMMMMMMMU���UUR�O��U��MR����������U��R��O����U�Ɖ����Ȩ���������訨�
��������
������






����������������iiiiiiim��������

���������V�NѣF�!B��Ҥ @���������N�`ӱ��l=��/A�+��44444444XXXX4XXX�z=�G���44444444�l;��c��R�x�@�CO��5؊�y��Bŀ^�OG��k�5��jDz=]�����iiIIIiiiiIJ���"""�""#����k��*����=qh��2�ok@]KF�j2�ɾ�L����X�RN�I/7�W��pJ.�䚲~�� g�%%��n�"�"7_|ܒ��R�ލ��R���+�r@v����������gm�a�wU���.J�$Xw���@�2����JXέZ�9��Zb������I�����������񑪲rZ�����������Z[{{{r	�Z��*******+{zZ��[{z��{rY�A15AA�UuuuuuuuuAAAuAAAAAAAAuAAAuuuuuuuuAAAAAAAA��������AAAAAAAAuuuAAAA;D��4B��Q"D�&L�f5w�'P�|fWWcTx�6
]������������������������������c�YH��4�sR, -l=�@+�kx��̤`Y��w=����.����k�$)�2,Z�t�.��T�K���aac`�����������IIIH��y��Iթ��I�u�9�7�
�3+�6L���REǬ~��� 3D���&#�c�cC�6�l��܈��;Pc�}�"�Ց�����
����q�@����paXg!r�%�J���LA8A_���I �gD���}�}�g��4c/6v�.����h�����v�	R����!ʠ ��$���++*������������(%����"��"��������������///////.�073���7+3�5�=�($���(7.�1+.�57&�000000000000000777777770000000000000000////////////////.����������������///.��(&����hѢ(N�*$I2dɪ$3$I2d�>1���F]����i��,,,,,,,,,,,,,,,,,,,,,,,,,v;�O���X�r�F�-���� ���d�%x��
�w=/e� jŠ ���� 01��)nl��&��]�������c��ZZZZZZZZZR����RZ�������Τ����=�t��cy�Z��y��*�kY<3q84>8bb28II8>kl���#X���7��ϱ$l�0�IӰ9��]��D	~�$7�hӐ�گ�xr
�f�7�xr�����>��%��u������IK�P}�u���(�tp���֏�֗�D)R��|��WSl� ��$��  ������������������/((/&�/&�/.���/00000000777777770&��3�����T�TF���ۗ�ۗW���^�ښ�����������������������SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSXSSX��������Bt�R�D�$�2	�L��2�t���+Ա��-r� B������������������������������c���x����a�����,l��.W�ij��	��-D-,x�^ޅ!!Nj�G�j��Ͳ(�Z�l 6�����e�ZZZZZZZZZZR��RZZ�������Τ����� %kF0)�q���s�{x�*�kVA0�1$�� $��7�<���E���R��$��$���_�OE����&���܂�Y��A_�ބ~�%�@+�$pJ�$R��Ԡ�$x6�]��ѫ0�IA�gd��׫�5)_�9!$Y��Z$����T��ͬ��0�Y ͉�$��� ��YYUUUU���AAAuuuuuuuuթ55����������������������������������U�R��<( 1 ��=�����=�����9������������������������55555553��������55555555555555555555555555555553��577775555*T��"I�$�2!*M�2	#!0��İh���v6K�����������(��ʈ�)g^PnDr�;^ޠB��-���1�%�4�v<^/�W`{��9�%5��-r�;�K����Q��c�����l�[-��e��-)RR)-l����""=�������=� �������	���h��+V1>.$��*�+�$�.��݂ϊ����U�U*Q_t���S��R��j��H�T�oaJ	Q�%Ģf�pxhx�pR��)pF�K�h��F���}��W�c�w���4h�$�Qa�I�d9։�L[S����O��PMU�R�����QQTWW���SSSSSSS\�[����Y��]Y��^���������������Y�ښ���	jƆ��JOe.j��n����JJJJJJJJJJJJJJJNnnnnnnnn��������ooooooooooooooooooooooooooooooooooooooonnoon��������J�L�2bI�&@��5w���et�wH�ӕ��z<^/�ѰZXXX444�,,,,,,,,,,,,,,,,,v;��B��ñ��s`EP`nl6�]�š�@xs`4 �X�z8]�ή��`c{��2Z�,z���<@-��`hi��l�[-��e��l�[%�%%%%��4DDDG77�v�vv��w6uT�����TUq��dt�4с���Y������n�PX�li,*�*�_:g ё��䢿�n����u��D�;RD�pk
��F�y"$�}�P9����(7�F��
.۫'�g�����/��:�j�+Z�� �$�07��������.���//000&��775555:��������=�5:����������)"""""""""")))))")))9�������ݳ��
��e����H��IIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIII�����쨑"I�&L�2d||Wf|fS"x������ǣ���x�����������������������������c��y�,�sz;��\�QMC�.P�W
��I)��X $���v6[-���a�G�4�E�r(R Z�x:��)���F��W+���r�\�V�d������)RRDDsssjggjjggjs{jM^PEo]Eo]nnPV��GF^����y��Z����� �>��A���U|`I,/x"�
��(%,9� ��K�6_�A������o���v�iv�i�"n��1����qmq���\ox= � �|B�*�����O�N�RO���WW��[�����������]]^������������Q]\ԑ��]]^��T�JJJJJJJJJJJJT��JKJT��X���Ĳ���Kڂ�s�Ka��-RRRRRRRRRRRRRRRRR--------))))))))))))))))))))))))))))))))))))))))))))))))--)))RRRssss*T��$ɓ&L�����f"�OWb����,x����aaaac��4�,,,,,,,,,,,,,,,,,,,,,,,v;�^��N�r#d��y@ᬱ�4(�u<gt��)�6�N�ca��p��
���®W��R�gU'V�J��k�9K���l�\�W+���r�[%�%%��+d�I����՝���U�I5y���u5��y�]�ek#�AJ@	&�*�i,J
�#}�(���Y����7C���`|U�H� @�HoCr�ǒ��H����9ȻSr��;@�H�_q�\��\��M��Fn��E����m.Q}���30�c7yI�4� U9U�	kbbIVU5KKVPjnMMnnjgggguuu{{{ssssDDDRRRRRRRRRRr��)�[%�nnnh�-��IIiiiiiiiike�ZZZZZ�l�KKK\�������#dh%�����R�l9\�W)iIIiiiiiiiiiiiike��l�[-��e��l�[-��IIIIIIIIiiiiiiiiIIIIIIIIIIIIIIIIiiiiiiiiiiiiIIIJ�����"D�L�2d���B�!#N���`��cб�4XX�r�]�CCCCE������������������������CN�ak�� 44��v9��W��oG(C��Ip��E�����.�
 M��*�����ssoRgg-g`s 	x�\�W+���r�\������˕�ZR��戈�������Zܬ�ԈΊ���Լ���.����ѓ�f�$����%�I��XB�/2 ��l#�+<�j.&n����a�GC������7�#}���������mD��<(�m�_�%~�x��O���1"�F�t&5�
Q�+������Qh�>906���%UST֤V�EV榦vwWWWWWW74DDDDDE%"���%%%%%%%!��e��v;
JJJE���`����������r�\�VÕ��l�\���`��snz:���F�^-��j��Ke��l�\�W+���r�\�W+���l�[.W+���r�\�W+��RRRRRRRRZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�l�������)))&LI2d�+�1����@��CCE�CCCCCCCCCCCCCCCOG����z=�CCCCCCCE����������E�����
e�����x�[-L��V�k���x���]�@�w)ka� � ,	w�)
�����X����#��Y��nl�/6��n�����I��l6KK[%��%%%%.nnonnonmE�-�	�Nl������hEY�UZ�X� M_t��܁:@��+�����-f���&�X5�4��"�o� ��;K���}ڒ ��1�J�Z؎�%�o$W�����J
��.&��	��߳*�� � %���%������58]]Mnnnjjggguu{{{{ssssDDRR))l�[-��e��l�[-��Ғ��"�Õ� Z���v9\�V�a��-nMsv��K���!c���l�\��CN�+`�$Q���-ggg	v9\�Wc���v;��c���v;��c���v;�+���l6��a��l6��a��l6��a��l6��a��r�\�W+���r�\�W+���l6��a��l�[-�d�>&$K�;���, z;�CCCCCCCCCCCCCCCCCE��������CCCCCCCE����������������O&�ȳ`%��z 9���;�CCK���LO0��ǈc�1��n"X�t�Z��Q�#6�ۛ�$�,�ފ�ԈR�RX�x�07������V˕��l�KKJJQ�]]T��[�Y��Y����bCV�>�n�s�����C��s�T������Ɔ�`���KzSt���	"伫�n���}� �$��qQLkJ�d��܍)a�
P�	a�)I�fjx��Z����p c���`���V��u�yy�������������IIIH������l�[-��e��r�\�V�d��,r�T��Ƌ��c��X�Dus)-uRz6^�.�`ӱ��)l=�CCE��sr!K`i��l;��c���v;��c���v;��c���v;��c���v;��c���v;���a��l6�+���r�\�V�a��l6�+���*T���CӐW������),,v;����������������������������������ǣ���z=�G����z=�Fȣe-y�ZR���y���!�₃�oA��J I@���Թ� 4��+����ax]ޤ怊�Z(X�Ml)6 ��G**�kR�������v6W+���l�����)))6��K\ۗ^�����Y����C ^�i՝4����$��P�>�KN�PE����J"���x��������P��}�ro�����Hٵ%���r!7&����(^E���$]-��SW+�d�XB����
�B�bq�Tۗ�Yڙ�^�������JJJJKK[-�˕��r�\�W+���l;����cŰZ��� z;�G+���i���R�� v9��<K/Gc�����z 8C՛Wac��4XXX4XXXXXXXX44444444�z=�G�a`�������������������������������ӱ��v;��c���v;��c���v;��ca��l*T��8�sı��v;��CN��a��,,,,,,,,,,,,,,,,z=�G����z=�G����z=�G����z���K^���J�o@��i���95��.�}�N^�nР�V���!� ���,--j5`-Dl���OF�%'�`c��H���x�F�/������c���l6-��d�����--l��0+)�������#F�@�| zJFb���y� ;��M����MX��[��[S�� oJ/����~>�����Ⱦ�Û���%TJ����B��"7^E9	 ���-I%��Y���d����p�b&C�Z�vC�Ȭon�nnh��jE%%%����e��r�\��ñ��v;��ca��,,z=�.W��`��` 1��,x�^��G����-l=-�a̱� XX �l = �UW]�MA��c���x�^�G����z=�G����z= /G����z1���=]����+��4X4�l6��������������������������ǋ���x�^/����x�^/����x�^/@�`��M�40�Uk2nl<� *�Ç*�`��R��^su` n���.�E�,副0����+�,]��^g2x�ݍ�+e��z<\ Bǣ���,,,v6��a��l6]K[nm�+k�Z��pb�&HѣFL�=��
)8fF��	�.ꂘ��j.���UX�5 �X��"�Xf�_�$A�"K�7��J ��$�/���0�Q0(9 �$IAU"p�6NV#:�pj��
.(:5�V��`��5IH�IH���l�[��a��v;�CE�������CCCE�G����r�8E����ǣİ9��  M{Rv6^.�	`г��� x�\ �f"�')�� �             �x�^/����x��B��ǋ���x�^/����x�^/����x�^/����x�^/����z=�G����z=�G����z=�B����!���`�`ӱ��l;��`�c���z=�G����z=�G����z=�G����x�^/��� � x�         =F�A �^�W*�a��EVx�=BU�ƀ�J*h�j�� QE#4 �+�� D�X�,)T^gz�<K]��Eg�c��X �p�^� ���z=�CCCCCCCN�'c��I���l������:�q0�Vʰ���  ���{�����X�4lň�h���V�"UB1d���
°�85�J]��L0V3R� ޿�_�E(F�!$&��ݥȟy�L����d�d���[�����Z2PEuju)))-----r��`������aac���z=�G����x�^�B���w��4�x� =  �!��"���N����	z��^�����rj�0QH��001��p�\.��        �x�^�G�ac�� � p�8@ �� � p�8@  �� � x�^/����x�^/����x�^/�����l�.�+����x�F�����ǋ���z=�G����z=�G����x�^/��       ��p�\.���p�\.�����w��=^����eTP�k�X�!�R�2Pup��M�F�(�a���E1pp��21� ��T���`�Y��^sl�[�`��HpHs�� �p�@  /��������᧋��i�l�X Լ�LJA��\F�zJ���c|,}��[�ׂ�3"���A
�*.� AJ ������܈����oa]����w)J\������)W����/�r6r&�v.�8_�*�������v<�#:�iՀ��mL��e��l�[-�`����aaac���x�^/����x�^. �`ӱ�� z�@�.���+�$X0�Ģ� �Z�l;a��G`p�p`p�aK ph`qJJ�pppppppp```````c���p�\.c���    p�\.���p�\.���            ,z<^/B���ǈ ���,,z<@�G����z=�G����z=                .���p�\.���p�[�C �A�o�E#Q�@���=�"�Sz;^ ��,�a�-��t���ps�d ��r���z��&�;ޡŁ�h-�bQ�����,, �p�8\   G����z=�.W+�QHAa"�M�(zB���W%ATz���� =ʼ�pj|p����
�q�ʖ��>7a�0:i��¹%���Y�����I��� ��U$o�+��0�Ԑ��!7IB7.�R nEwV�-oE^unr�^o7�Dt�^
��L荗+���r�\�����ǣ���z=/           ��ı��l��.�����			w=��0�`e�h�]��z=CE���b� ���s�,8$$$$$$$$88888889��p�\.�$88080000000000000000000000000000000000000000001��p�\.�       ��p�^/����z=�G����x�^/����x�@        .���p�8C!�������������������ǋ��,�^Ul=E�@F�@^�w�B�!h+��,��,�p��+���EW�I_�����CJ篦b�+�0iʂ�	J\�����X�%��y���7����p�^.�  ��l; ���c`�H�*�b�'/��0 �sp(�ҫd�Y�A�ͼ���J�
� ��.d�H+��F���]�HF�$��ą(�~;Vv�� �Hn$_��%�����r7i}����� �F��ӶM[��� a���x��3��6����ce��z=�G��  �X�z<\!��!�����%��� p�Fb��`s���z9^�
N��ȁ'�`P`!��w

 9F������̒�,,,,,,,,,,,�z�BE��BBBBBBBBC�C�C�C�C�C�C�C�C�C�C�C���������������������������������                                BBBBBBBBBBBBBBB^���B�B�` HK� 4XdX T8��ެ
(.�,l7�H9 t�]'B��A�Ӳ
sPR{@q{(0�����XX.(0 4Z���y��!!!�c���   x�^���c� ��\���=cWBȨ㧝z�dȍ Q���ƣDTUWQ�c���K^H���eW*��ХT�йEE�D���t/��(�F���(�J��0h5��d���݆帱A��r"���֤�(IHB�kGhɓս�-��r�  8]�����x�8\  ���``ppppps��� 	g]w
=E����`K���	 	w"7;���^�!��C a�s`D��Ey�4���,lQ���E��������������7s�XY��z�=E�����������������������������������!!!!!!!!�����������������������p�\.���p�\.���p�\!�����������������������������������������7�ӛd8	��x
��� ]!��qp��P��4� � ��4I�(
���]�1@`�@1ux5�
F(�1?t�:�;���N.U�@(��PX 88���y��z��8\.c�i�4�E-:r65�Q�N� "��'=*�(���q8{{Msl�-fx��8�	o7O�����܅����_�"�$�����ӑ����,+�)E�]�܍�%�W�!y�}�jo���7aDi5��;۪)j��K�;���*�Q��5H�5���r��/�   ��� 	z��C��!���"�Wp c�I���y�C�]�W��(�y���KB] 
O���0�z=A�������A�G�s�խ�0�w;��竹��w;���s��,�y�ޢ�W����z�^�W����z�^�W����z�^�W����z�^�W�����������������HHHHHHHHHHHHHHHHppps�0000000000000000000000088888888$$$$$$$$X$X$X$XY��z�^�W����z�^�W����	 w��� ����]#"�O1g��e-��,WN�,Z2������t���WC[{�9��{s-/jM	t�K����p�`ca���y�����!!������@��Ǡ�k�����*ƈ�ѕ"BP$�t�X�r�FR�{5]M{)RNtwV�����%�a���}�/��T��\�(�$��.�(�1 ��7������0�+��U��F�
�Yk��i����:5�9�"�)3�9�"58^/�0080X8 XP%�,�		z���0���c�\ X%��z�Q �@����.����g�K���)��w<�ޮU��w�#�hh8�dt�Y��y��o7����y��o7����y�<ޢ��G����y��o7s���w;���s���w;���s���w;������z�^�W����z�^�Qaaaaaaaaaaaaaaa`����������������������������aaaaaaag����z�^�Ws���w;���s���w;������y��o7�s��0�y��<��FB@^ A�0��`81��y���EF�QFUA@ �����*�#?,`m3uv"*�
���-��^, y�<�n�s�XX$$$889� �	)E2x�w=���Z�q1 kP�-�I j��"�5���6Z�d9cP��!j`$�j�,��5����\E~/���]�"�%
P%���}ġr ܻ@@^H7.�7�_�^HoBn	BH����X�HFUu4�ͰX�R�.�q�4���5V�`HK�$�u� � 			w 8E�.�aag��P`PQ�.,�z�<މ�ǈ�����$X5�.�w�5�.�=��ÃCF������qw��e�4�x1/�����������������b���g��\PPPPPPPQ��y��o7����y��o7����y��o7����y��o7����w;���s���z�^�W����z�^�W����z�E������W����z�^�W����z�^�W����z�^�W����w;���s���y��o7����y��o7����������c��000.,�t���=�Aޡ���  ���dc�W�(P������
1X^DXjڠ,0�,)	z���m�NQ�p����P$9�,�y��o7���,,�,z
���@�@A�d��q*� �  B�E�"����SE׫�4	��*H
d�  OW*T�/��}ӑ�K���a/"���(��M�P�t�t��JI$lIv�v�a��H�e�b�Q_�梁K��YƋ�%��Ơ՗�ӬBXp�� ,�x��6���@ 竹�� -z�]����Aqqqw���.�y��b�CRѠ�@ �!��a`(k���6ARx
<�ሎ���{��0.,�4-w=E����������o7����y��o7����y��o7����y����s���w;���s���w;���s���w;���s���w;���s�PPPPPPPPPPPPPPPPPPPPPPPP\\\\\\\\a�� t�������@�!�Q��a@�� C�a�.Ԁ~u� Q�r�S��FD��],o��@�q�� '��A{�,=U�1�ܠ��w�� ��^n瘸����w;��W������c�1��]sl($�?~�q��$n�L=���)ic�-�k�P`cp:C�(��*f$Da�c1�`\�P(�J �k!$��d���l�a��K�Xw�7Ҕ������}*��M� C`��;:�K���h)b5��Z4�z�J[* 	�Q�� �p���,  ��w=^�1p !@�H`������\%��x�B^��@C���*+�%�1-�PM w��6[/ǘ@(Ph���h(;��1�.000000.�z���������������������������







<�o7����y��o7����y��o7����w;���s���w;���s���w;���s���y��o7���������������������������������H�K�5��x���� ]�၀���c�h(4���5Uw'cWHWz�NH�dD�{�ƦJ*Z�x�)$���R�N����� ����z����瘣���w=^�"���A��K����,s~����D��)�U!M�J����r[pK����e��(α���� �I"�����ӑ��Ð�I!_���O��_t�wv�@$@Jt������A$wJ��X��K+N���=]�n�W��Ս�Fu���y�E^饋��/1qGs���URw�
��^-��1��z;��� N�xh��xa��zR���,(,��,
w����c �CMo1a�  �����  �  ���� !wp��a�0000000000000000000000000000000000000000((((((((((((((((((((((((�y��b����������������������������������������� C�x`Se�U�(怒�(�x�< �K���$�3����`C��`4I{飤�QPQ�JJ���Sr��[")%�!a�`%�@�s����sM)v=T�#�W��������x�<ŀ  ln���/�,Xt匼����D�Z�O����P�W�����B�]&�{� ���}��n@_��F�(���xn�	�9��P;I�a+�7wi7N�A7NDoF����O�J��\R�\��큳[;é%��J3�߀�@��BY�Þ�s���y�

����h����AA`�WH@ �d-�"0�v ��9�C�� �E�'��P�D�a!������P9�00�x�
=^�OP����{���w����{���	w��!Ws����D(	�
�uw�:F!�K�$(,(�@�0�Vf2U!U0���D��n��08(ғ���9)z8S\����(�-L�� �gphk�A�....((�w<\�W7K�	K��B�91~�tsа�&�)H@H�"Bv�-�7H8@�Q�9�P���_ḗ�����n�$ ��oc{�@+�/�@���q��v%P�������H	@H�nﾔ��0��+�����I��.,&:6[PC���w=]�Gp�ĥA��y�

���<ۛ�!͐�{�tX4\09��w����9^� ��@���W���;yc�̸%���0�Z�r��:B� �]᎑P�Gs��
�w�:C]��{���w����{���w��������������������������CCFCCCCCCC@�������� ��������� ����������������CCCCC@���@�CCCCK# �L�Ia��"�PG��4`P(��{z� �BNQ ��:B���
b����R���۞!
��"=	w���.�.�`෩EtE� Z�

w��59� ����o1����,�v3�]�N�'�4�֏����QQ���r2P��q���pQc��,���t�D 	�^�a_t�$��iB�.��.D�NB�_pn���_���h�*PrW��0΃2�1�rF�gآ`��	-�ͫ�O0�Ƨ�՝��}�Q��A��]�"� N��c�PPPP\\\a�R����0�x��o1G0��Т�(+���)�4�)-
l�/( ;� C	�I����0�!`כ�!�.(�

w���;���{���w����{���w����xhhhhhhhhhhhhhhhhhhhhhh��������������������hhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhk���w��CC]��{���
Dcp�>
����ΗHC�XX<0,X<e�""(��1=,t�������N��`�����י`�$���@��  +�PaA�Mw=���r��e�0e��z�<�/��W�:�GG~9��(9�����6Rx���8E�T���H��FW	_	�SvL�K��T[T]��p�.���Z
��	���l\��8#b��PJ���k����1U1x�e���MD	EMZ���$������Hk�%�,...000.(0�v"3�;�F N�P !qwW�p�`K:k�Ҡ`Z
�2gl�<
]RA����@#��ף�=�
"�?|
w��@���P�W����x<����x<K���t� �����������������@C���w����{���w����xhhhhhhhhhhhhhhhhhh����hhhhhhhhhhhhhhhk���w����{���w����{���w����{���w����{���x:^ ����(\d��2�e�FJ�t�;�� oP���  ����2�6�a�)��@�E�� �.p���<�*��ޢ헙��s�r#R�#��
 ���p�5������F
]����  !�x@ Kհ�|=%h��֌��~���+�}<ܡ왕^c� �w��c��`�r^
F*�n�������NBo��iB�/��&�(��1"�����n	@H�7&�(���0��$h��@��n]���r1��.B�/*��p��9��AU%dOd���(<]��,	y�=F ��CC]/0���Ap@P!�WH���v�9W@"�/��*��,��z��/+��Ss�!�Ԯ0"*�t�n���2�HHp�+��(�t�B���@C���x<����t�^�@@@@@@@@@@@@@@C���w����{���w����{���w�;����{���w����{���w���C���x��<@ �Qw���̦UP<4(d< 4�� #y��;
��T�*G4��2 o�t+Y,y����]䢡O� 2�����THSv 6\����!aw�R�:h��-��`��
y���xh�	���bz��$��:��7�~�z�\��Sf ~�)w
);�C�K�ԈD��d�v��n����R�$���J	RH��4(9/(1�p'��g��B!}�gm�v��."|o9��SF�$e�����`�.�xCe���w���x�hK��X�(h@@�� ��8�X)ʊ�~
�l4��2
�n3^L$QXܧɎ�QWxphXP�(s�\	��WT1"x��;�A]! ������������@��������@�N�K���t�]!N�K���t�].�����x<����x:Ba����x<����x<�K���t�].�K���t�]! �����t�AC�FC���R1x�+�4�
2�
Tx
�����*g*��d�2L=W9 x�<I�t��/7H���<i�i��{Ug)z�ށ��OFuV˥�F�l���<�{��0�x�6T����4,�֬d����9�̰4i�4RX�F�A^19*���g%Sώ
,F�������0QQyX`a$��(�HW�o��E�����Fo	B��Sw��}Ǒ/3�
;�B�A�7�����b���Ԥ�x�����N���9U5�
�w
"<CU[�T��B�H������CN�����kZ)ՆJI%��q�+� pQb� ����H@�A�(Y�x8(�`X+�(()��t�B��������AB���.�K���x<����x<K���t�]/����x<���ǃ���x<����x<����x<����x<K���t�].�K���t�].�������x<C�].�P�wР)k�<eQ�J�x� �������Q�*^M���C�e��'��)�{�9S����O���g''!���B� � 1v�G��F�P XղԼ�4�x<��G�(�S�KX�?fh>�:u��H�/��7K͜ ���w��;����c��U��E_��7��7Ҁ��&�HM�ܛ�@�� F�#p��7�D�ݠ�A�}Ӵ� &�oN�}��Ij����J���6�wz��0�X(<�Ej������ m�H���C�P�{���
w����^�@���OUd������ވ,*�ov7:� 9@^�Eˮē5�����)t�6]IIr�;�����Gx{� ��D<%���












t�].�K���t�.�K���t�].�K���t�^����x< ]B�!N��HS�)��
t�����@��H��^��Q`3�4�'�8��T-]��p��X�E������doC��yx9� ZA4,�F�L�����!�"�7����)R2��� �@�� !O ��#3���`j����.RZ,,..�usr\���kDlwI�֬d�qW	������Psp��;U�I'�b��%�N)K�PJ�. ��aXgl6.��,0��v�*T��Wĕ�I_8�
����$��0(��]��hÀ��|v�,Z�X�T��� ��HaK`e�"J�p�;�
WB�] � � .�'�U|�d,��"�n@w����AE���r
4�-VIz�;Ɲ���c�@"�P���jK��R�	 P	9j{/W%t��3���>��FFFD@B�  ��!���@@@@@@@P׀@����
�t�].�HPPP(((PPPPPS���t� ����������������������������������������������:C�FAB�� a ���G�x�S�TP04��"
z����@�LH�S���+=��� $�W�Et�A��¯0&2��n��9J	ib!�xB�[;YK`<(��<	 �-0�Y-��,�z;��E�\�� �@W���.ެ��
����G�֬uA�I���p���g�
��2����C'����X�b

�A���K
ûe�E|�;o)@����h|`6(�΂�%�_(��I,(�7��ð�$AaA���%�H��(�D�/��쑿Z�r�z��"��UcPE�GH��P\�%��v<�DF^ �+8sR+�)uI��w:^�7
�p�k`����z8\*I"��P$@Qgq����D-g=w�>ǌ��ң��h���nR"-m}� � �wK��"
00�ka�
F�E���@GH+���t� ����� ����].�H((((((((��
*^�/t��^���B',d�͇��,\����e�;��h�izu��Zu\�]�vO��ׁx���1W��c���^�rZZ���/z��<ؑ�(K�� 1�0�9%	Et�́p��Qg6�À00tg�C��2�����A$OQ`�g�����s��n=}:EDA�[�#a����a�$x7�p7�r'h��HoF�oF�7����Y ��ob@7��Ӵ�)E�7&䐹�>���>����Qnz�BB�]/d��߿�^~��Z�^r�7
�"��!�P� qx 8@8 8;�`���l~�Vz����L��@0�B50��EWC�(D��F"�uMMsL�;�Do3��Pp'��и��%�{9t�H���a��!K�DD=�F0�d\Ew�^N��(P((P((( ((((   ((((((((                                       #�<,( T�P�dY��Ա,Ѽ%�U5�2D�.(**�/"R^h�f| �QٟDD�V����;�P�z�������dɌ���o'a+�X�\P�5��l��;����7�7�@�8xPP+���sl���9E�Y�u�_�^r�r��P��r.�y�6����qP����³�D-�����A_���^D܈,+
����h����]��aXT��8,*R3mt��i�좖��t8��՜؁�^����ѿF��*��N�jow+d ��(����m�*�m���Vt�w�xX((��+�P��]�4(��R,0*�2K<JQU[�ݎ�&�*[dd�H$Y�.�`-,w�����!C$A�����������������A�{Ũհ
..






"
�x��������I%�x��<� #@!.���.�����x�w<A�^��	���D�&�T<d�:�S�7�u��1���1z:QBG?"jP{ R)x����=K�E ��!�[��
0��
t������$�1wC��+:>��2@�C����1�й����XX�=y���B��U3�	'Ɍ;�_(��8� ���7��1$�� �&10*�J.+�m���:Pci�ʿ�����Xq���;�h��^���w�K��׉+�B�����@�GQ���w��A)��8`,�"�V,-	w"8X�S�CR�$Р���I��,�����{j{qy[�@����M�з6�G�ѝ�0�	r���:@C�H�@���@D@�KE�_DC �����������#�<]5%���z������ �����������������������������������������������������������NN@]�񓗃�1̰TQ�$ ĕ����,�1Ml����;�<�E �V!=?|S/S%h�Lr��X"�!jj�E�m�×�˫S�����4�
R�uz��������+��0W��<��r�����"�;�r�_��h�UT���T�&��`�)Jk��
%�֨~JJ��ؠQ;d���K�7Cu(^H7q0��>�~�������v�@�����/��K�_��l;	7�	�����tnA7h�]������]�@�`�v���#�1"}��aB͆�[�<(0��(
�.
J"(�w����;�4�UE���4@//1l�[�N���ÄIX�[�U�ޡ�n�UF3Ћa�P(8 D8�4�E�*�""-l:EH�BFFFFFFFDDDDC�DDFf �k��b �� �b!���"""""""!������P�@�@�񑑑���������������������������������������W� r ��Y�x	�0q�9����jbDz�ٞB��],'XFF	O�DA�>��>�S�F��8eb�+3{1��X��`]��mUn^l��)=[�/ѡq�c�I�5��U���XX�x
��=\.��U&�|�
��-�0��^,�G*��ܤ���^r�ss"z�].����]���_g�B��ȍ��� +�%�/��D��n�A���$$"$/�nI�7swr#wJ,%���M�QrA���}��7_pB�À1�4��4�����	@�^�O�A�x@�#���w:D^%�i��A⠃E ��wTU�'WR�Pk��f����x�,+�X,�5���Uؤ����ޠR�@6EH:"��� Pv=.�B!P0Qgac;��y�0�
y�����������������������CUZ��^�p0�������@׀���x ����������������������������������������������������8X��ӰPD	�
�~�
#gnEz�:C�g��Q�� ӑpV�W����Д*a�M����H�����uq�c�S�0A�!CАS�� �׉xs��J*bJ�z������+x�8��pH���480��i����r7�3$lo�֝Y�F�H
����J�$�!y�E]NJ�F^z�(b��I_%.*o�"�]��P(�[M���1$������L2E^V>6<Am@>_8����&8���(�����'d����Bc�����8EECA Cj��@pG�P�):"(���-�JWJX�WӋZ)�a�4*�v�BA\&G����&�/b.�b�oe��4���X�Z�.��<p�� & /��p�QP��R3�0P�pppppppq�������HX�;��P<)�Y��w����������_@o�0@0��q@�1P7��,dDddddddddddddddU��%�S��r�ѳp��]B����K����Ö3�#F�"H*rFFAc&�ē:���%%l���&��CȞ���S�P'q077��A|��`�(Y�
*R0
�z8K]X[+��/�#���w��2d��I��,�  �	�Zl�:@��`hh�uBVȂ�(A��
$�A��%�$]�ؑp\�;d�ȯ�DoyW�	!J�����_��(�.%�K��a�ڍ�;�Qq.2���R�ք������a����S`4��,"r*�p������2,z*�x��@E��TS���w4֣�k	r���QVȈ��ܤ�XIK  ��L �ҦD�"��x�䛦����$��dVvӽ���^w��������>���G/ �j�! ��@�� ��n�@���Ơ&��"�B��n�B�0C���e�
DF2D22�x�����6B��H�FAB�B�����H�A�B� ��� � ������������������ � !C*gY4|W&L�d�������1h�F��SUE2�`��3��!=/THTSfB�91ق��@�� ���s�b"50��s����v ���6]�1�g���dj�j�x��J�x���ȁ�	+���Ǜ��7�9���bu��2w��ӓc
{Rw��^�o0�ѐG0r� �A���F���NB��JR���A��n���Ȅ��_�~�J�7�W�H� $�_��_�W�oF��.����v�%�$^W��$�"	7&�A�0��/�eqB��[�i�30 ��)��	w�*�6R��	��S=}:���WʯT�W��K{�Շ5u7�q�ѡ7��xr�s�y��Ɯ�0��Ј�P��@8���_�/$WP!��2���i�*.
r^�z������������C!�aC/ W�x�ɸ��R�9?	 w����@�/�P@W�PI�`=��g}�������������������>������������������������Ȁ��H�US})�fy�Nz@��D@������ B��)ִW} �������B�E�F	K�HƃB	IFB�N�B��0C� �A�tɜ4\	�R��0 ��
=	
19x��B�CF��.�Q���Y�ձ�X;�h�X�����)�,<���2*�9��dF*b�9p�/���pr7�7/��.Fn��n�7+�r�r67�h9����"�.B�)B +�J#_��0�B���/��Pa���6aXJ�7ܑ�Do��z���7?=�kBo���hX(���..�w �>�F�@�FH (��=[S[,@�7a�S�,��a4�� Q��iY��̈��J������a��r�z���͑B'ә�{�!�5��
?T"%K 9w�)>�^�i�p�P����8 �h�x���\=I4i�(���,`�T��,(�4�,,��#"t��������������] �o��XXXXXXXXXXXXXXXXXXXXXXXY���+��P��Q�d�F3�&�4�@�F�U�����
#v�������Hh�kD(H���NTɧ}3!1=}����^a!��W����i��p��Ս��0��b$A�B��@7��D��<d�%��v���\f~�=�Q��4*��r�K�09�� ,Y�*� h����{�<	,��h���ހ�d�������������R�-{`2VK8jRbgD){nju{^ojuK8oo`@A8U@>L]8r��� ���V�2GF�9S�#��H#�9y���^uD]Sz��;�O��]��N�p�8�e�U	^w������=[  M�PS�[��dļ%E��MP����t�Q��D(���8^ ���nUP��Q��A�˪�ĥ��^JR!v6�o��Gx{��2r4D~,�SD,UVx����X�B�A��@�C^7y�(��{ Hw�=LNA��IA��FH�O��C�=�rJ*********DDD*r��r����\� � ��K�:�-��*���Hs�H��U7�2@ Z���_L[�ΎƨT��\��Up�g+8 bh����Ĵ�$i�*Z��,=Iz;�J]���qPq@� ��AW��U₿�ƄV1����d�F���K� UT��	T�	TSf9%M0K0Qkqq3_<�KʕJ��5�8��RPO�J�}��d���`����a��E����a.E�I�)��`E� �6��F9ի�OAF���Wx�D��� "b�#%/D<n)5z��C��ל���E��*�̰e��.2p��&��#K�dtd���<�;0�{�$h ��m8|& 0�%w�)���/e-�x#�1� � `HH �
z�����R��1PS�!GV� P2����p�?	 t�����CF��UL��lr�
S?#"w
����=@NOH�EEEEEEEEEEEEEEEEEEEEEEEH�EIIEBȈ�Bȕ�R�8�	FH1�/"1ht,T\�a��bp
O�Y�2Tt����=}1�*U�Q!����Td�!�2֏� �ӹ�*0�H:"bF�z;����ȍ�doB�a���l����������@C#A��!��!X^��=$�_%
r�;EB�T����Z�Uɟ��� (�>�P0��n���}���(��B �,8�o��H��rW��yR�t�)BoIB����Ro��jR!(�fA(�]���aq�{�T d� (�8�_��KG�H�K�FX���CB@LC^ ���y�{�1��J�-U8	5IVEx�����.�+����6�/E@�X�E�|��I>{&~��Y��w���cMŎ�F˥�.r��  ��x(������T0Q�l�X22F("J2��%y�*�"56BB�H�F��B����.bb.�p���;��/�jk���=?w������] �礮��a���}>�O�Ы��DD�%""SH?/w>��$T:*�ch^A��Rd��:r�#cc~@I7�gJ�$!SS?9 r�LJ��+��(Y�D]�j��1B�Aw��2 Sз{�i�܀Qz�]C�A�d�!`C �����N�/|NUr���d�a3���Vv˹��S|//=gW?9#"8Au��	�$�av��R�n��Ȱ�%�$&䐾�Qv�%���0o}�"v��;I!a.��.L}�c}�p\�p1�yJ&�h��u'a���z�X:6���k�@��N��XY-HDEUu���R2�.���?1#l8CK�۶�D.b`sl�����>��]!  NV�3����"ެ�$��8#�� ���iA�0���L,#y�������A\/0�@U��S�(ї��8�x���,P`us&^%���A��z�g 9x�6	H���)���@���1W{��J"2"�)t�����������������
�������EK�ȝ� C�4Z�M�8�KR��,leZ��_OV� ���8 �+�+G§N�Z���t-��B��ޤMů��00���P8�色0�9|W"W��4�	 y�5� 
;�.�W�x{�e�(�qb�b7��:�������,b� .���H�O�"EP�����TF2df`�b<_PU��\I.'���	m�ƥ�����ͪ�ʦ�)(���#%cV��CC�#��"7�dD�`�������AV2 q%�4/6˕ʀ����{,r�������LDQ�E�)��/g��@$����(�-z���("3�9T�X��]��%算�����l����8NY�N������� �G�V��b���.4��.�WWt��C"�%�/S�WI{��L��!��JM�8$4����"	"}� C��KNT�BA�C ��PwyIH�`�Ōd����#%#%%%%%%%%%%%%%%%%}
�>��H�H�OȈ�	���$>��>, U��1S�n����2-�E���/P�0B���OPq�s��g*�'&^"rJ"�,h��P5jP1%h�#/d�Ęhp�hAh�ˤ,,0䔍�4RJ������HC��`�F�$��=\�� � �ߐ}�B�x�W~��<]5(� :	$���QQ.@U5E^gMMsnVV000�+��+�A7�rE�W�[jU��/�����%����t��,HCS�KJ�-���@$k�ʞ���K]\����,Ų0�22��JZ��v=\.�0�@� ��c�+���bow�<݁a�  ����k� E�����T�E\A��(���c?w��A�QOSAĂ���*�AE�Ɓ���'�f /0 �pP�s�`8�����?%E`%T/"//1=1%t�;��_N��'x� ���D�<�]�^2Dr
(XZ�,T1})�����������������������������������<,"#T/?Z����G�C�LLFX�AǤj�@�c!l�O�CDS���UCV2S*M!Q\�3�As��S�B��0U��S������2`w3��X�-z�3�NH��/��˩�����_G*�`�&���ߣ�d��
���"��Z24�)j�O_OGl�0�|oyD�k�R���d�C�IQI@5VkyXs|oa/�HW�Q}�t7XE���_�&�ڈ,+��I�
�F�E���HP����4�Te��H��G�h2�,,���fuD"x�D^��7��u��R�Z�w�
�1��^$@訯7� c��*��l176[Ug�� 9R�N�0G	K�`����g-|
f? J
r�w<Nc���0&�c���{z"�����:��X��%Ep6����D��$K�+錂�9������DJ*",
"�%?TS �/};�"���"'�g�A��.�ҙ(�)))))))(Yy(x ��x���B���OP�Z9e'� �Ep��7{r'`#Bj�	ܡd��^g'!A	G/�δ*�U��L�`U8ˤ(�E�5�Ĉ��]\P,d����@+�A4��"� x���6�ֿZF"���N�7���'|c9�\�`�Q]c�"LOβN�9��ʕXa�o�\�������r%��;T��&&6������y�7/����n���iDAr3zr4�n���^Eڹ ���~;W�́T�و�55�ux�` �ُٔS�h�K�$Q5�z�	
p� �*�v(:��=���C�B�W�a���`����J#�	�5�!UnPz��6kS��=�O�����F�"�r�(k�$-��^JAPQ�X,
X�pd���}>���CJ��1AB�&�H�Z+�P0K��TT,���ML�4� <�,��p��NFEȌXހ!���H ;�E��"//cw>���H�����������������INIA�U���'Wc|=TWcTc| ��0���=�F��l�N�:�zd�����^^r�|r�X��U	�r0ut�����D��/ @��^�$���"$D���2��/W����D\�a�y�E*� ѧ���ݑ�P�{���W8�ѿG~�;��2��x9�A5��| �̱sKeY�*�"k�|PpR��Ъj�l�f�/��S͌��O�K���T�T��X���Y�)i��OFʐs����H` *�<z���� ����\� A�n�0T+8��x���P�.�*(�44��v ��� ���)j���h#��� l������*<\� M
�T# Px��R� F�e4�a�M��S���((�d�$���%��"1f&2�SW%n]y��^�ʀ�����(�`k���bJ^0 �ST#cy�;� �i�%�F�z�����IC�����551S��jh��x+�- ���������������䌕�FF�// $��~���^^���L��fEV�j�(J����1����Z� ' z�D��\����r�T�B�I
�M���� YX�SH��#�%,aL��,
�d�X�|���h�"�*����5��"X;-7���'&���Jb�ƅ��P�X��ք��Qpטh#�4e�"0�t�\.��[� ���0 PY��y�K�@@W�J^	&��&�J��ŏg
�(���E׫�5�v�<w�Y4 ��o��]���n1`���w���"/��3�>���JY�]�x��) pW�x�y�Bk�Q��u�h-����4.�h.��2��0IpF����O52P�ЋRh��P�Q� ���09JEaP���C��8$8`49��g4jz0;�!o AC�dd�"�6�h`� x��c�X	��rALP� Td��4�
�v
�����W�H�DB���NNNNNNNNK���������H��I]!.�1'��g�LǠ�DG���?F�q�;�ѿLĩASP1�"��C��Wc*Е�F@ꘪ����NFE@H�C�S���B�!o�� ���5ފ�y�; ��[���e%6`s д/�a����Hެ
O1R`"t7�ѿG~�9�5v7�f*����f:��o��f ))��d�V�C4�g�(����Z��a��Cc����༮ۀ�\�bH5�pZ�J.�2�U��Ģ�3j`<�9�,�)��#�&�Ƶ�:u��`PG�G�(��<d�" �=}�)�������B�Ġ���^�$d����Q@�W+�!`�Z��c��Z4�c:(�884 ?}"�OC��ގ��0�A�(��ï��	��v<�G�.�7�hQ{����v ;�	h���H1�
� ь,P����,Q�X�p44�b�2jv*�>��B�H�R���Q@ ���P �p��9��20z̦rrrrrrrr^^^^^^^^^rJrb^*��HW919x��������W:U"ɣDiɃ����W=�9&���5��� alm�+�&^rru�Ӫ᥂�"�j������k`	`"����Qi�����.�A8A8r��e.�ӳ���7�:Oɜ���u�ѿG~�:�s�ve5w�K�Ν&Ʀbb��dpQ(���|�yW��x��]�m*I(F�;�û`�%�p#c�A%*pg6��(0��2Z��d�)]os,l�"<�.-�~T�x�#��5��sp���%��P�wҡ�(h��P �X�#ʒ
�E{%z��]B� ��!AM� '��-��"�,^2z����Ӑ:��Q�R�9]p�=R���"��9���&&5��R��C�cyhS���2r��Ȟ�p
�kqq��JY�D�Q�X
JA8�rP24��0�p׀aI��������<T���x�3���L0]�T	�R�T�UP�dd����������������ļ������P� � ,�BB��xZć���ѧF�H�Qѵ+���# zb̰w�0��gd� ��S%X�r4+
�S
bv�#/�S+�`��1�,��E��Tt����) *
;n���4rPrb��)Э*U7���':��J�QM
u��o����Ɋ:�	�c�d��ny\���D���	"o�a�7���!J)K
�R�
�cb��!Qm(�E���R�0��@��1�R��I`J[j
��h���hꇨO^d�"����$�o�� 1p00��S%�F7��+���`D��x���K�P04)��Ly�5����T�IC��^
�'Kނ���@�N��ǫ�I�_������:�^�y����@�S@�Ac,dE���QK�`���w��ۚ�Z����A\����ljddD�$����ЄF���@���j�����"' .Q@�a�������c|"w<��T��OLOLNH�H��LH�NLLK�NK�O��K��K�U��C�$��C�2 �\T��-�TJ���y2g%H ��dz������Ӑ~��˔-�5%,8\\���b��*��=�JF��b��h�<u/m@>wx<B�������o��*�X:߿F�vK�*��94�4�2"���K�nA�-j-��� �p�v���������0���J�$Fϳ���b��U�-uIIA ������������g&D(��l)�'~:15��b�d��^.W������\ ePEx\���HT}�������*Nk���h`1޺ZR�N~�RUz�#r��6���G"�.�"!�` a���""=5v�ٚ=ޡ`��G��AdOR��]�h��I�ە���%1"}>�E^�E@�Y����G���e\�P�@x�h`*�q��(�@Y�x��0]4T�%8����

Db^bFD(�n,ouz
;���@e�jg�%��&%�o�&5E555C��������*������)�9"C�Ӭo�#��Y���H`y���b��d��X�PD�JG+Z���%�<PšS�� ���2~�w6��I��������LLL@P ->8_>�#+eL�0h<���,�Ӫ�tk��~���,B�����L�(�]�M�,�T*�Չؖx���ުX2��@]M^mmQqt(�+6��X����RM[�RPX�
WX�B\.U���%�d�R�����Ҥ�x�,~,
��(�f&��8E�D�x�B���4�8� ����Ub_(�������9@�����%�E��Y��՜��U������\���#�OɎɌ,)��XD��g m4t��Ŋ� `�o ��ǡK�=�4b��r�����
����� :[&!@!�Sc��׋��2�A�H�wЋ;��DX5���w�������O�F�^��C& �����˹��z9SO/�3������55EC2R�4��3��5553�����54�uw�AɊ�0Zv���/ɡX�M�{%r7Hs����@5rbU�= ���FG�l��].���S�P0(�5��%|&�#|}1��<��Ӄ�"+�T0yT�W�^a%����b�#��!~�b7�~���!N�	!@�4���p�y��t]y$��%�Û�)@ܛ�
���W��IDo_���M�	}���M�5�_Ą�aDD��  �Ɇ����R�i�K�ڨ�uD]��It=\��uňɑ��!*�~�z�r�=x�Sw�������� �B�{p[ ��vB/Q�a���j��5UxU������{<Uz;�A�$��:�Fz2~AP)��M)%-?*��l*�"( �;�MN"� F"T��Ƒ	� *@o��Ca�E@�Gҹ�8����ȸj��*C���0Y��xh�p#轌�� ,JJ""
J�r��l�)"<B�H�����ONIH�LU�����OOOU_@ag*��'��g*ij��j�H��-P}k!Ѵd�IvH���+R�w�N� �D���VI�#SH 
?y��$��.�H���H  {10p�x�{{� !9�T=��Pt\��~�5s	9@r���c%�D�*;��ߎ�b�N���,%?"/ x�*��J�-e�D��yW��H�VnXH�o���~;SrHXK�%	!yR�畅a� �/��\��ƴWacڱ������M���Ph˔0�ek��ѩ�*	H=HF�t� �=DH��y(�9h��y�"
.�v
�9^�����E��0ǋ��W��xq��`l���t]�h]A��E��J"�x4N$H�a'_[!""��h��%��d����Qr Q�n���	܈6@l<��adi�\��@��23�W����;�P` I+�9��x���f/ ]Ur��Tg^1=H��4,�ST/??T|Tgx�)��������**W=}�+��W1%#1""?cTcH11cfc:r^L���*�����Q�d�]P��b4*�ѱ�>�R>�Љ?:��� K��!i�Aŉ��
7�(qD��Mr���)�}��>���+��?P~�0,.����uw>����B$I�߿F�vK>3	*��rF�?z���x(<E� �$B�(�I%��a�ӑ����}�iv��J)D������t��}�W��r4�7Ct��D��&��n���m�}��m�8+�t�+��~��ph	�I���'��ɫ�d�2^
0"�x�����#�a`�;�T-��XX��---u�,��8x���Xa�ϲ�H��k���X�$�Z�l����!}3-BM��8`�Ɋ��x(j�9k�D\���;0����0�w((��*���1���$ ��0����19IU��Ӭ|#z�<�.PS�0W``#��yl��J��!ʚ�#�Xh$d�QL���}�^a��$��NN@�Ȉ�O��]��F�`��rzzrrz�*�9=THcc=Wc9#TH9c�
tKDv��N%"��7��uGK��P��b��d	�*!:L��E�o��m�AEX�Ixek1( )x͌uA,�C��B�z����|9l�������\� o�ݐ얿��o�d��MP���e���Ȉ*���Y��gj�XI�rx7xJto���Ȱ��� ˴tn���w7q��_|�/����})a�E�v��s��*�0���ȸ�����B~溤�f�p ���:w��¯�g/� ���9x�����1u9:�(�(�20�T9ul�=�DEה!��&�g�O�W��K�_N���g��bױ��2��V�5��)�#w��Y����y���������� �.��A���)�(��Ps{��\�%� (�좪�|d�u���d@�  @�x��[�T�K�H5��Xl~D�F�^
(�#Pj
,g Tc9w����3>>1����O����X�P���B�bH>3��������
�
�4::4gG*��;J4hѿ*rD~bM�{��b���]���h�ّ�&�bz@���M�� }3,ND�9&�t�S�D�1�*����@�,D��� ��,�i��1&��d�
�߿F�vK��Ў@d]�XX9�@�f�n�0w���H�sб���( �"w�����7{� (<,�D(DD�
�9y����N��`�sڳsY�;`9�D��8ꄧ)P�1/x9��&8OH��OWHk����w �����D��ŃާeU�r��1�b�'�!�
��x���6 �B �9J���F�NT�E����]�g��ȓ���}'z9��//f/H
E2Vz �������I�����C�ܢ�7���:�I����U!��В��sכ���DU��^̦rD"�#	%p�5������^݁/Qg�@Y��y@!*C��2g ���b����
jj�eN���*��K���e$֧d;*ԄhP�e&�i�4l�N�N��1VB�eY�ʾ32}?S?|"	x>�7�'f/w����H�IR���A�,=p���������1px���qv� Z�׀"��C��a���jlc�~���9?N����S1)�$g��f&�+a����,v7��*���ȎR�U�U��STSV&��H�֪�l�`�t:�\،K�W�"
ciA�1y���z��2��XљM����Н}�;�CR�]%�7aبz��W �"z$�x�$�:�	ZM 1z8R����o��	�1{�4�!�x�JU	��y{D$�N�sd�^

�brt��0� z� 
�X8��|�v$x�5�T%M@%^8"]aK�^�_�Д�]9���z��y����֐"F4�W"9}����'� �!BW��[�aҦX�"%/|%p�����*|WS=Sf&^D�@䕙����A,�n���Zt���Z;!З�>�:u��X����UħZ��Q]k$�7�S�&��A�;���	�����Q*�/��E H�I^ahU��.�AA�RҊ���y�	��Q�t(�����!��'ą��>?~�1�,c&��3�G��$nTG�c2��@�0���TD-�H� ��T�6$��$�J]���Ѽ�}��F�� ���)F��J"��!v�M����L5P]>6gK4Ds>2UE6@>w��16��zvK�ӣ&Luv5�ē#=Qh�z�9Q!̀ 0!rQ����ar�J	��(	��=9HS|AyM�!/mNP��p��(X�dh��ף�<�D�"	d^T�����d $D�w��� 䚠k�X,T]��b��c?p�&5�5�8��8��ch��Dz�"NM���~~X�"=T(�����^c�����d�l��FBl��U�� Hh$�]����t����g�
�����g�	���f&TK��9���zb�M��#�#w�N%
u��B��%G�Y�2ϋ�B���Js����iߧ .�1S*A\d�;�a@�
`��`e���d�!�J	��a��@!��E-�3����Db���
��ĬZ8�RTه~���-|*�9�%P��<E��B�CSO��TJ)H��#{�I$\�>��}ڻW�*��I��R�� ��I�>�	ݪ�rL�y!r[T\�Br\���Iq��]u-t�J+���j(^=k�ŋ�֗���\���Fb1�o�y�He4)��t�<ށN��c���m)ooj&r~2�l
���@F���D$B�e �H�+ŲzLD!�b�d��TN8[���a)z��A�'^o3����'P���N$��9*�w�PAxPY�E��  �F��S&�dTG�$�L��a�jwq�dY�(Dƨ(�Z
�f�w�� _AC ��!�Qf��(@����`��"t�"��!�ŃBΑң�2�����*>H*L��2��X�$_JꃐN�i7�,�EH%d���x�( ),�ѲX���3�,�Z@�aܮ^u�w�դo�������
;�Kȉ[�$C,��^+�''�n�-���/3�քE�ǲN��v�_���-Nb^z�@�F����ʺ��%�1Yyʤ��ڠ�`��J�J�"ܻRE����J/���tn����u�^D�܉���n����Ⱦ�Q�	!J.�(�K���P��q�pF�n��k��@�Y�ڹ,N�R�p��m�	NA������ЬrZ�Dl��z��]������Ry� )( ��� ��"Ł���nSB���F�zJMIp���xd��L����X�J2Mc���I�x>��:���<4(�L�M:@XPc����A!��x6T��Z� -�X�2"���U����l�����T���ou3�G{�TT40��\8)�0XZ
�)v9F����Hh ���� t���� �����$J��ąv3�2�l����Y-:Ъ@�Hh��_�&ё�fa/ѩ��/W&�G��G�Sw�%�$1
&���B6�aP 'K�����3�IP�шa+�	{X�b��]c3��,��,�*��v�J�Z���;%��H9#?Wfcfr�����NƲJ��7��q��;Wjo�\ ���a�7R���ӑ������/��nB�)@���DoyD,8޿�Pc�o�ĥ�JA�m��A*�6���L�P\�]\/�Ӭ�&LK���VcT/#Tz���:B�[-B�$9C�ś�X#E����{	a�@�����*A�Ѥ��V920cB�oIl��S�?:�S �
*b9�V7����Pu6C���T??TTT&����a@���X�@Qj�ȳ�ʚ���j��v��BM��e�L�=��<�P�@4��Qp��9����������J�/7{�1�Y٨ �=��9}�KJ�/
w=BB�_F'���31�*$��3����d"T�A�Z)��?cB���0*u�߭tu�i�#~~.22b�tu�V,Nt�����X4 ���MM ���B�E��#/�aC*��U��Z<�B� ���@��߾��DBЃ���*:Ӥ����X��C2gH)�� �=\!.W�˫``	�t�����l��&���k��*N�@s�4Q�0(.�"%x=\# ���s�Q��հ�S-QRr��"&�6A�O���%�S�B� ������K�s���s"1HN2���l%�����ˁ�% �g'!��aB���Ӑw*!A��^K}�$@j�^� V�HPpkԛ�QP�s����iQľ��S�= �t�]\q�4Z���;#���93ђlb�!����%UgT�Wx!c�Q8�S�h���%�a�ak�\]��.R�M?gz�Z���OG���Frr
(0�Rx��^nU'Tph��X�P�(X%�*rƮ������@�1�γ1����	ZM���wèR���ɂ�c"/T},F������+������:ttk�*ѣB"7HI��P��H�2QQg`����P1ө�����w����E����@wTW{25����$$N8�ߎ�js��BY��/���T#�����#t�� �;�E�Ŕ�ƀ�������sqiJ������g]g->>k0q.>4^oKbkI]P4p
�A���U��g	Rmg#h�`��ĕfNѓ#6f`pP4���ȔDG���h`[�*l��z3�6K��g�N��8<�,���J����^�*�S��I�)(Ù�h B�+�� �p���Z��Z��X��U��,	:ë3)��)���:�zAc$��	�4y�
6Y��.�-F�
M�s���,�"�jm�	|S:L4��R^��"y��@n�aA�V3���������Z�T��"��T�'
�H�x9xS�X�*��H�$��ɾ$&�&~@����B��N��~%jq�Y���ĳ>�dUa�|t�_C�Н&�jw�㎰I�[PS�I �X��b�j�� !��ӬT}���/@�p�4@Ҡ @c��h[�qIJ!��lo���߿XЩV�_����-kA)�N���'���K舱��HQ��30�a�yZ�M����
Qq$"n��<��v�%ڈ+��m+��v����Dlf��-gn]U{v:�"<C�*%��j �#S���FD��hʁ��)�ʨ*M]��9"%v >=\���&����x�����% w����^����U`��^������h�{����y�2(z0ukE�'���E�������?w��� M;&��,b��-
� ��\�������'�x���7��9WT:��� ���F�r������3Awx�M ,�`81��4R�w���=����cxa��ˤ,T��dL�66b3>|H1WHw�)��h̐$��	��FHI_O��d:�FS�hǤ�F� �MP����ю�u�V,B�^*RM!�%� ��N~�u	:�u �I����D!�X*�4qAKgLVT
4l���h2� �=쇣j4hѣ�ňI�T�B5Dכ�dK��p��%%�ϲU�A�G|��Β�/�r7M�a	!}��A_��Av�04o$]�K�䯝K�a���ΣM��F��j���%�`�)uv&��ѿfeZ���2¨�*�*ƨ20�Wx������26w�<J@Xԗ�'��b" / 7� (8� !xx��ŝ� Tv�H�	����{?*,2�,Uyub�C���VX��1��ؽ\�������$��P����U��E�O��Wz����f|Wt��*$+��,,�:Տ�@ά*.�"�rJ$-�
0�Z���x��`#��!��!ȳ����� 
/c/
x��&�vD��_�����!���xi��(c������*u�e!jr�Qٕ'B$I4���H�F�:6D�eLR���ߑ�>2y�B^���B�rb��㯠G��5uED'.�+���0s`5�� �ԜeyM�8�F5z��ߧB�:=��*#���J�5Dt��ےD-e-��Q(
'Ĕ��fHXK��/��RM��%t�	,)" ����	����4IJ�A�������	�Z���Y�Ôآ��x��MJ]��`�ȟO��d���*�GZ��դ4/y�#B�/�DAA�"\��V�P�`#�(-�XF�=z�[� ЉfcySו_���D��6ϝ^�	�V�M!�#�)�cj8=|/W:*.�X��9�{8"Ar�jd�M�ʼڑ^� ��	�9)�S`���A1߿NF���
�ДH�x��+���(�z6�Ρ
r�T�g�c��2'�t�0��� �%�z��w�:H� �2.L�qc��л��4�P���&%�t�ѣZ�bt+Y,:��C0��*�D�_
��_��߱��9w�dJ.zT��qΌ�;�`'�Ф�BbD�@E���
s0_$8OIN����Hӌ=G|c&�`��2F��V�V�ѣ~;#�*�J��F�|X�U{{>>RPJ�/�,9"��/��H��� ��ȍﱹJ�H���,$���ܒK�,I�M�`��rx}Ӑ��t6a��ț�ܾ�ڸ��PE�_Ag�TTV BR�5���r�u]�
v��2B�%�뼁{�4%]����v*=������ ��$�	)(�Q!)�#��t������v�c��H��ag'/�3�������$<�u�����,&���E,X����6b��ꏧĀ�G�ɂ��D������
AD^c�e_B��o����%��2#��:���,�,
� 4�����p�8]��秣#/�WIb#�(���P�Dd�D40d��zL��BAlg��!Oz��uff00�eR�
?&Uc�d:1�4N�9ӫO�&^*�H r~�tk���i��U��2==:t�1[�8,�t�Σw��$�;��'r��9�JBCF�N���!�R�	*��*����	:��F��%��|NtD�( 45� �55-|�F�d k�;l+�0��Ґi!}���;k���.�1�y]	K	7ҩQ� �%��R`.v��Lؓ[�U��+�N�c�N9xC����.�|&A�:��H*1�Z�b1ΝB�2DJ�p��S-9
MV(Z�]]# Wz��E����a4��3�a��ǰ -�C��� �	)����@�� �xc钺���ʤ3+�Sh�d�u�j���J���ɘ�����!�m��L�ŀ�1SՇ,gX�H+��-���Z$4\`4��B"�^%z3�<CݎP�נ���$T�=��z�����l8NY�H��|ScH| ���2��,*zrzL���@	3��_���	B�:4c�Y�9W:����_J�	��*�T�4U
�#�?T�&��5�?
d�\I����S��WciH|4<e�Xr��`bPj>v��c��E�ŏ��N��z���֡N��4hѣ~�`�H-*
�jz=_C!�"���h���x@������(^rz��zz�t ,ļ� �BκK߿�.
"0

�,x�
��F�c$���^�OEG)c̈��Ѯ-XT���%�Q�Nt��+հ2zJt����52P����ɩ����w����=F
��@�Ɍ�C���B_	Y�P���r��sx���;��UӬ�GEI�% daM�D�Z�t�H�dtP�vbb�Us�@�'a�#�)��%/t���َ�������Ӓ�=="?sH
t��:]�����ǡHа��ɉhc� 1�"�1T&�y�;�H���D^��W�Η�:zb^L�7��M��d�~��JthֲNb;$�Vt�)ӧH9f*���2�f
/�b�jb�Q�;:�ɒ�@���A����	D�1��AC��E�	%���Q�֤� b�[����"���@0 �����ɝB�%��ѣF��-dЛ��������y��F^���S�YuYuU-�H�hX`���v;W�д��R�MuF���3��E,`�f֕M�"I�F�@J���R��+:~~tu��iRg�`b�.�50vdjȋ�E��ۉ��pGx�ސ*�w;�_J��/PRPՉ�)�����E �mH��O �E""R�+������UA(�Є0 �I�Z;�Ĵ;���d�32��,��ERP�rQP�5s�&�`��Y:�Hɪ��*��U�*��<Mr����=Q��DO�Ƒ�Nfi-�W�;�P���: ��s���{��0�t����
����:��J~�MPvffHĞ�F�'���br"�����1R&fd�r
�h֎��fF��!п�
�@�(p��dΉ ��v57�HS0���	��g,p����C�]�0���s��E�և��Z��QU�߿\\\~�7�Z��\�D]�"J.
�r�>�U���˭mg	-ȭ��h��-�W��}����X���U�
DJ�#"Sp�F2E^^EE`jjb5%TZ�k�$A*��bDt�l���'�ŋS�&��
F�*2b�w�"�as���A��p�����@�CWp((��i�Q((X�`��y�50�&62�G� �����@�J�ā� X�B�;F�Y,H}������1�$'|?B���F*�0bu�� ���P�@T�� ���Fr�z���)����U� ���e����Ǚk��(�	x 9^����s�a�J�=w�<ȏH���	H��.�p�����/�j��gI�Nu:֊b��ѿ�#G���;��q)��N�:uv1ѕ|f|X�	�w�ߎ�S&��"y�� D�TS=Hw=�3�\�a`S���.""��
}�>�`�h�SNu�uE6EY_���ߣF��ũѲ&�~*�B^*�l6]�n���AsQD��-�x������
z��[�\���"�ǋ�����.��l�j�� �ނjZ�o463kl
���}�&�"9����Z@��L�#Z�jӯ���b�AI��j�GXT�h�(�f�z+=���^a�g� �"���4/����W��4,� �.z���Eq)m�/�K������!	Ӵhz�%�q�1�!d;B1��(�$�7�G9|NFr~*�%M���H�=h�
s0V� P���c��FzzF��ғ�d�������W=l:B�dj��-��Wpz�ʸ�������P:������4��S�c1WT&9hy)Q,eX�4|X%�h�N�N%��h�Z�Iʙ)��
�|d�:u�ٖ?��s�c�FF,~�D�#}/"�����7)����9��C��^���W4����K�� (iV��$DAf$ɤ#=c?tx�,h��4o�,Zuju��~����2J0!@h�$^� �U�%c��f��V�p�����ޠX�	z6WCF�i(��)��e�eQ��I�p�j|\�w����r�D��]'/���Yh̞�`��V��K��kհ$����Q)�C#��n�7���:���ù�b4�11 rJ
(z�D�H�X�h��A]��AH)�S`}<��$��$��&ɣC��>
� r���"��/UA��P��V2=9WTX�,(<<��\��pqf��R���hb(�	w��FFC]�� B�g/���E0%�qv'�R �1�c aa�x@s�<��<�������"�X��,%�b$��
�4 *J4@��Q$�'F���KY?h@�님�#~$�!����ǲ:ub6g��1�	1Td;E���'%����9+�1�*D^�f&"Xl(�6-RuE 
R~�0��b�@�B@�[�l̟�*����w�ߎ�jw�ߎ;&L����ľ��0*��=r���N�W�$�Å���1|���A")g	w<CC��i)c �}Y4ռ��f��z��Æ�Rt6��ڪ�ּ��m[�]����ю<t�O�NA7y�(���0x��$�`�N\! #N����ကoW�b�@�QWШ @)�=�
�(�
F~0"Jts�p
�7��QFBUs�&��	���D(�Z�I6EHвZ%���,g��!�r����D�B�	��d�}
��>+���D z��IS�-SS?�,�l�? gr��*AM�
�~0�f|T%y���Ȝ���EIE]�P1Wx�s��<]�̮uP,�ro�a�%�Z!&�D2F%��ɋ2*��gH+�Z��4to�w��ߓ/d�c$o�dA����Tc|�<M���. 2�
�"w���!�o+��.�DPgunx�
;�ƊS]�����7���Y�*�kZ�� w�ѣ~:ů߿q�2w�hT�� @�W�I)3�{:�yĢ�qt\����Zk��yA̤����Ԋd`��ܼx�}���PT��`g���n��B�"�e�!�XX��}�~�:Lw�Ѳ+N�;��C��'!,j��aK�u=|bVz<�b���S��)�¢��%.���ʸ���5s�J���&�SSoRup]�&@aeI�NM�1�$�ֲ !�Ʊ�9�K��!c&7xC�Y�:����%&F�,1=-|F�~z�b��0�PQi�P(H�@��4$�DAB��`�df ��G�!� !gp����fHx�
�56"�� ���IDO��NI�cS ����Hw��Z%���$' u4(Z-d�qsX�r���b�3����F�\���3pt�� ��	���{�\dT�e�b� r4R�DPw����Yܠ��i .��hs�c�U��:�F�W:4z7�~�����4o�-N�
���y�#�!��E�$����
p��n����(��#���w���A��
����	,)%|=%SWT �D�/T&b�	w�FN@X�h٘ǭN��6��1Z���,�ʡ�+��L41�`a���,B�.QWx``���2��q/���4�WĀ��J�)�����*ɐ��( ˸8�)U| 
F;'�ѿcy�BC����P�&�U����C�c3�m�&��#=/%w��^�6��@k�� ĩ��(x:*�DD��U�P�PG`Y�P� �]�p�,�x s s{HNT�,����	
x���������hU��2X���){A�'X:ţ�HcN�������HR	f�50p�R�F�Q]>:uuq�@�NY�	�|?N�PH���S���H��@�X����C�/PFˤe�~�Ht�H�
�pǘ@(R�'����?d�����oѣ~�q�7��5ì�)���-aW��q�XT��YȚA��/��h�2r�*"(�w=CFA^�����"��6(���̍��]�T׫�� 
�9w����2�d�!������E��@�K��l���2Z���Dgv;��'�e�i�FP�=�)����LO�4"*�/W1�XXLY��s Sfz�3?~�b4bH,d���s�Gd��$��h8�gU���=h��Js���k�Č	�^M�z�L��A�(xi��	�AT�Hs���|����
9^ƛ��"���Ag�I��H�K�B� D@���B��_D��D�X;$�V�*$IRhV;$$�,cu�S�\�Z���ԂR��ɓF���L�1Ѭh����ǿY9
t��@�Y�B��/1S}�����H�ޯV�rXý����	t���
= �JT��
��@ �b4'�v6C�F���F�7�8�ѿ~����"c JJ
�Ԡ�y��=T ������N�e`Qc�aԤi��l���Z��(�@A<v"7��(76DKτ/+����d�a��f����x8#��i�.Ur����ǬZɍ
4dAΗ�H���x���I�F�XT)͝��
/%9?"=c1z
����Y� ��x"
���>�9EɄ���C���ȉ_�:���T��5��ь����Xu 䈚�2
�B�,eY	/&:��0Uq��C��0�p�Q"���G���b����L<���8xȖgp;���Rn`l<��ט�i��wH��j��c b�����R5655s�?hu�"
�Z��F��Nɒҭ
�XL��������m���	N�:�hЧF>U5��>�� �ѴNA��l�X�^zƐ~r�i��jy���&9��
��6C@������ȅ��5C�6a-�*�q�~��hѿ��hѣF�4���#[����3���7���K[ם�N�ǘr �b+8������E�>{u2{z�=�
�����Ԡjj�`�k.$���A7�)�S�X)��gD?hzu�C���YX��CF�������B���@bc�j�����z�
#B�� 4��-Ld����r��w���'IJMLDi��%h�d�DH�������ȋ֬���C�V?�7�A�$�>��_EO���GZ�*��L�da�(�b�F�Z�  -���04��D�)Q
�����(8˚
Z*�(�D	�b�F2J"��u:��0�2l�iʊ���2(V�:������Z4h�9ӨS�6�Ӳh��;�F�4o�Gju��N:֚�-�~L��ǩ
b"��""Y���:t��'V��]!��.�7���c����,}1��#%
z������ �fd�iR�2d�w��F������!&��T4����ӱ��ܝ� �/ �l$��(<C"���
J�N�T�%��c��p�p���z������ɫ���6"KZ���*��:�J&��I
P6�=�E"�­3&���ưH�G�dDF,l�b����+�����	�҈H�!{��bz�bF"D�P�D��TQ��@�]�"�=M,H&�/9H "jp��33����*?*�
2n�'�9�e2��v��,}�;0�� ;�����0q���xhXs��5w��U�� LgY�C@��ٙ�':���A,Ģ���,3���!�2~D�})���$SB�bª`����ŞI,ZM�ň��d�����������B���ߕX��:A�%��F̄tl�>>�(Ѿ#BrTJu���Sf�==iF�~2���9(:��r�3�c�1���A�P�Ң�梪�7����H[��8�dQ���=B^�a7Ř�2~��ѣF���;Fc�R��¤B͓��7�hx#�+���K�j�:Z#�iX��|�;v�J���ar)aJZ[�r�&0 ׫��޼X��8��\XQ��7F�n�a\�n������,�i̽	S��l`ढ��iH���Г:����P����f�Uf�)���=9,Eh^�r�T��Fr,~z;��x#�(9�ɡ�@�3�Vʣ�xJC�U�-3�3=`��b4dٖ�d��V���k�hUbq 23Մ�������Hz� z�`��m�C �ZHcTh$�	蠉x@�h!*�+�4,E���^tJB֋�:_Dg�T1S?Z%�r�ll�,�Y��:T�3�VL�'h�:t��#F��ʓӾ!�Y&�<�"��$LN�F��u]�1$�VtT��MjB�֋LC��'1l�(;���H+�A��J�*^.�
cct�����Z�
��,aՃ�ѣ�!߿G�ΝFT`ը�(�$�ܕm�(�%�*�	تھ$�,)��r�!��J���;k��HWゕ5x��^Ý�No�3;aꦪ௒�Ė���T "�;a�%m;E�_���Nz�m�ec��H���ǯc�k��D!���]nz��P�RI�����Oي�9=:b�c|}d��(C�\�
qξ�ʤ4Ww6C�Χ!�W~� P�6L���F:5����� B��,bY�r��bt�;���?1t�����Z4/x �NЉ�Pqb��n�C�'6d��LIU�Aɩ��h��ɒ7���b�
��>��gK�ʝZ:7쓭h�:Ӫ磲X�:t�Q�8�ɓC�ʳ#�Wi��+�h�;�� g�P����ED��NU�3GӼ�9erl��|
Tt���
h(�r4�w����z�9[  J�	�B��q�5��-X�:�OѣF�u�2dɓ&�,X�����hl((�2ul�V�g���z��w�� ���ޢ̈́����JU�ל����UC�T�A�h��=*���X��Ӷ\���Q�f|YWS~�
Ɖ�	�N�������@"���x�:�NAH����d���E��C��4�y��#@�a@���s�+
���H�HOOGh�^^�L����bT/�J[��oѭ" �	��j`R����I�����$* 73��I� �~"�����~rr������y��)���
�����N��� P�lmȂ�DG& zF0�X��UPdE����XL�"jm�N~*~�a�l��N�@�A߿�"��F:ֈGd�jիVQ��2�w��e��"�#�S*���r�о>����Nɒq�D�\Ѫ��fT:2d���KȔ�ɘ��������;���@H���������$JiV�d�d��&���c!ߎ;*���4ułD�|S*@�2kV�,��%ur����A@��f�Aqv��DGrK���y4�f��\!&�M��Ґ&�Z
�7� �B�ʿ|cv*��P�Q���Z�*��t����l�֕z�ĭ9�ý�^�w��7����������<F	�+�J����lb*�秦"�B�$g�$��e� @�s��1���Hz�F�b@�N���S|F��1'_�Z�u��	N�R�1x�$����FTUP�P�C�se�(��9=|9
	w�;�$jd�, z�<G?:J
�o&~rF"�t���W9u��H-:�Ш�ȁNP�Wh�
6BS�6M�N����q�X�j�L��G~�;�h֬F�K�6f4��_�Z���;!щ#ThU�u�d:�k@��0�4��~�L Ě�r ��"������;�(i�(�RRz������N�b7�У�HӭZ�c%�=�%��G~�E��PDU�x��� SW�)蓑��aHs��X�nD
#I8z�)3�[
��,M��7ъ����1��\��`�ZT1TX�ڊ.~���2
�Jb��}������&�z�:5�,�:V-F�G�ً���K� E�D�A�C^�D��!�����A�LN@F���I@�J�XШ�!BU\�r�'������c�XuA֫�F�1��#:b��j�)�bo��b �5C�caj��K����^�/���y���c��!�X��	�T84i���J�~��*��5%}�����	W?:tqߎ���I�2NF2~u�6�ֿd�j�zƍ��d�G�Ō�~��=�q4"V,[fX��>���v`5u�u2	� Ď�v�έ�X�L� �u]�4�ɘ���!:�"�"b0��h�,}8C��P�'�3�+��6��B��4�ӧZ�b���&�������F�4k_� �d2J�z"̅L���� 1w=F	U�^`�!B�a`�hp8��4�Q�X� w���" �;
Z��^/0W��ߋ9� ���?HWSB�PM	T�v3�`��VV�XM�@�6`��w���h��x�yIK�9�x���"t����9�"��B��-�W:�~��o��D���FƵ Mh�~M�����Y�#Z9�7���Z'*�b~�LJ@ ҁ5va �G�[3��"Ԛ�U ���Hw;SE�K ���MB#/�NAJ�w����< �T���!B��%5rY#�5�ʭN�4o�4B�h���6C�*���8�2~�7���2\GBMc�쟕&���ՋQ�_HYV��:��TZ<s�_֐F�e�,Ʀ̍
����G�ᄆG"��7Р��4"w�������C@�LY��b
�ю�h�֭N�:Ռ�!:$��2�PS�IAAAU��Τ4(
.�y�����Dg���J��9#S*:�xAK� �8[�<��հ�{KMjVb8`z���
A��3���u���!�`n��w+�F���
JA] JB�����!�*J^^���	3�"JʼDQ�"p�9\BLAU��.�AEqPusP����d (DD�)]�1+���:7��l`F4���[B����U�N��2�3�B�Bc�d���Z��B�H�̌���"4[��]�,�%�� ��0V�p��sd�h��Az�!��N��B
�le�b�!C%R
�:� H��{�&D4N����x�ZX�k'�ѿZ�u��F8����֬�N�F��q�	 A�2���+S�d@�c��rd�F�D���C�2h߲ I1�V3��`q�#e�T��\�8P{�5��}�<K[! AkV?~��A*�Y#`�X�;F�Y;%�S�B�Kx������c����A��j�t�QaM��N����LI�<-�`Б@Qw��-]�4L-¼��R���
,w0);� ��1�*'dL�ɉ�¤^�b�~�^b%8��"�P�h��-Q\M�Q*iT��a`A���_M�rHQ��,��ëp�X`��1�ȁ_DaDi
��S��������N8�ɤ�FL�a0r6f��f'� ~�i��ЭB%j7�I�B�����%�j�Z! %bà�CbU�^n�j��,??%tX�9 ���12 @G%��K�Y�~�l������I��AΞ�����)������*^�H�X㎴qӧZv�c!߬B��8���?߮.W(�i	P�z�|�;eX��R��'W"}���+�*н\vHӿFu���-k�zj����YQ�B� 0�
x<��YÆ"$c����ӎ�qюђ��-d�j���!B�k�W��F#J�aAB�CNWT��l�|�������fØ+$��<�Ş������Q���	�c:�K���X�v;�]["�ɦ���.�C�ф,i!�OԂ�6]!�`磮���bŋD�F�=M	TiĎAAq��`.�0�6�F KLF�UɁ4��p���~��T~�UP�J��b�,""�Cє�h����§Q�ZI��~��q�&��B�t����:8X�2r��hA
��F���֌�3���/�&g�Ka��  �%@�R�P��Hk�킇���*p����������%w�@Oٟ	u�T�c�bOQ�~<t��F�b1ӕ&@���ߣG�4o߿ѣ~;&I�/�#F����&�֓FT����'Л��j��� �����Q�Z�1/ѧF�8��(Tac0�Ѳ
�� �����\�x��������H�ѧ�ūV2���߿~��u�Ή����ƮL�k�PI1� �+���#}����=�)�%O��Wl�%�-y�4�ښ��꺘h���R����91z&�������[+��S��t�R(��MQ
�;��5Q�N�
�B�X���UiU��?Z�r �C�	T}�������*,Sp�=�-G��hYc�ܮM��W�bձWʒc�CDh�N����ߎ���U�X�~r��q�2dA���ūQ�H&z��- M <�-��:��(
�SX�K�t)i���b��`�zaq���
���8"��37��ҫcW*
�cX�L��:��&�{��o�V8�߿F�q�q�q����֬F�c��V?Z=�uCҫ�h���%�k_��HeY�-TcT9�8��H���Tf	#9K *���l�&��B�U�����������߿~������X�	Q(P�:$�2h�P0!p��p���%�(�-,=l6F���A������a��U�$��K��XDn������y_f�#P+ѝ������p��7$�"�����		z�3!z�&��N��"�L��f6er
��4W/cB��d�:�k�c:����?%&@%40d()����������¡`� g���6O�Ѭ*@���a�ή�j4eV�,����e�$Y��cC�,�Jb�_
�d�0,U�.bb(X�u��zF^�%��(�Wh~�.�x>�����K�P,U�2�К�2��N�E��|HW/}��d:6��g���ĉB��9R�#d�q߿~�jŌ����ֲ~������2A�kY?N>��:q'V���jՈT��ΐ:�~�
L�d�j5���%x!1x��%]MI��(�pQ7�;��,I������߿~���hѣF�4tc�N��U��4hu� D��� ,���#H
w�����oWxa�F�"){Ev=�[&��K���)gE�0���Qk4- p�[uu2PG���]IA�X�R�`kE	sAz�T9Wf~��et�d(�*@��rmX$�v�࢏0���$�w���N�����>�F]��#�#\\\\Z�U����2d�j$3��h]��Ѭ�?*�w�ߣ�N$��K2�Z!*uh�S�B���3�1#� l=�]�/��b#�g�b�B�@��j�# aAe�U;f�#{��2DD�Jƨ�f&�;A�3���XuLTŌ��p���ɼ�G�hM���K�c�~�4zի~�Z���닋���uG�HV�B��	�'�u��+V3>ɚ*r�!!iU�ʎ���b�WH�xHʸ(�2RPr�<N��6Da�@�Y�ӱ� �jŋ-Z�4hѣF�어Bu	ӨZW=dbL�4$X�P)�D@�2 0� �2�AVt���KJ)�GCA�qVr�K���KJ���7�7.������^NP��0qa��Q����ӇS�"סhp[s��gE*�r�ߓf~�����ƈN�&A�� Jrb�V�{��*z��@�P+�r0�+�A]-�.,��\~���dƸ��2S�1&WHt�%94c�N���j�1/���TпF��
s�ў��X̨Jr�,"2��l6w!fS"=Ml�>�FE].��+��D�SZD �J�SWf#w�&���O�U�&~X�t�<C_X9��S�b$�X�c���C�G�ѣF��d:�ZЫ$ku]��dF$���'O�4��T�kӉ�A�P��$�NO��CH�	z%"�s�#`�I '1�`���)ЧZ��%�S�F�4hѣ~;%��!&$�D�H1�:B�CF��� ���{�9��FZ�W6Df1K^z79^�p� @Xs�
`�-c@��-�P��dX$\]��,�����Pk0Pl�+( =�9����Ş�����Β	УF��952V7���dɕWc|B��)��-z��ӝN
zЪB��Q��q����니߿:�����5�ŇJ�eZ��XD�c�r"�|u���w�Z2���H�B@�:1'GW&�t�����!n�7��3�%�h�g`f@Ul6[���0�аs��0GyUr'�y�A��(8�������LS� �Ʈ�c:��z�H#W��q�XѢ���!%���h�F�4hѣ+���b}4hY':U
Ջ�h����������r	Ʉ�&�&̯*%jA�)(�cx���X�!��P׀s�$`� ��d	�̱������d����߿~����,Z�8��4:T�@8X8Px��{s�`��r��U���t��;����"� B�i&JJ��D�Cke�uͲ�x���ĺ�t����\!a��Ņ��ʬU%��T����+����2D9nEt��h���d�����ɾ>4F��5� K	F]�(Ъ?S?|*��
�.?~���k���������~�u���l�ߡZ��d��ŇLON�9Q',�Q���1�!N�
��о'Z�jՄ�IN��EN��RD{Hl������ ��A��_B����@���1QGy*�7�J�x��t���V�AM\��IqI�D��hV2X�|s�;��ѣG�N�c!ߣ�.Y4N�d};,q�I�'�i b��OOP�2���"�I��Ȫy65�o�A�pa�r�{Č��)��z�D_A�-��E�Y?G~�h�8�;��X�js��� �A�'TT�K0���8����D(,,J*b97H��Z�yX�]�T״�4���Y�5ռ�y���(Z��x�����(7�ޏG�Hb��j�������nRz6PXQ	@��
�����"N� ^����63�oѭ����&�{E����$�A�-��GY.,X���tu�����%����H�u������4j�Ь�~��Q,��HB�`�P�N:#�NU;��V#hF�S:FZ,J~�=%8 o����.��@��(X8��".b*��D�T����x([���N�@���F7ţ�h@�6fc��up@2��g)S�N�:Ō��X�c&C�=7��rbN�X�\Z��;-�4kG�F�w��V��đ>���?T|=#W|c~��~�U	9�fDDB�ޡ�E��A@������2S����Z�9֋cC��2dɓ&OߎɒūJ��S#Sz�n	l��%� �2Ї� ���Z�R ``�����ϳd���_+��M���&TP��d �9��ox�=>gEl<ު���-L���p�H 5�1����4(Gk'�K�4 u�Q�$kN�B��Z��f�2���]e�D�t����L�+��?�*�������F�9�v��0���hӝ&��$�H,TY��N��I�ĴX�c�ҥ_N�6������Dk�|X��1dE׃����6>"Lx�;�$�,*dΐhM\D���t��I^���lkc� F����B�l�_LN��Z�%1��.?~��;~M>���լ�ѓ9d��ՋG��!~��=�6Kk�FE�D�"W����P7щy*�Dg3�Boʳ1���d,M	)(! y3��Ā 4�te� ��ZX���-N�vKV,Z�KW�2�gN�H?|B�,�z��C"��@Şa���s�-�U�ֈ�t��5��	D��5uPgUb.t+<��HLڜ����E��NǨs���w�
=O^ƀ\͛M^7q{����y�	���g�Ȃ,dk�ʭZ�"���h;Bо3	N�j�0�3�4)
iΉ:����MakQ�DJ��F��GX�z������W%9f*=PJ�aSҤ*u�M�j���fiZ������_������6`����")EG�4�G��Q�7A��/D �a`r5%��R���J��1B�z��	cWY~T��ք֎�I22 �H���
�D�������/��4N$��hѣ?F����n=���D�ʓ MM�L�M���Q	��:u�դ��Ѿ;�Ğ��9
9h�DD45!�*�e�Q���Y?G�d�c%�
�X���$�>)���f

x3��:��2���Z��^jg5Q0.`z�^���ΪNS3�TF�#5q�c� �(�ceX�u@�|�1(=�5;����`�V���#��9�ʈj�|����*��jX�����Ą��,��N;"��&L�Ջ_�>�U�ɲfHc TJC��mC�n�M��H�@O��h����L��..#*�M��AP����KJ���N��;$�P�*;���������:�u
�3�@�@���Q�*@9�@H�P(C���.�"r��j5t��
e��!B�E� �Ja�bUF�Y��B�c��5�gYS9%"9SH=
��FH���Y?d����i�3>,�ӡdȩ�Q�X8��F���w���ѧWSH Tꢢ�ՈO���~�:����ٕŎU�ѣd�3��A��"�Z����o�#~�q�dɓ�K2XЪӕhT��s��lo7��i��w�b�ic��Q��I�(���lp�HBF(�`^D,o{6>oRR>t.��K�\/7r*��bj�i�{{��o�J\��op��ǘy��ù�Z��,l���=�">��%�\�@
j��ɤ��H?*�A�2ƇP�X�k�*�ɳ	��"Z��	���\�R+K�@���~�qptvI�\�L�*eN�eNtw��С`�$-B��ThTɉ::BBq$�㒒�*+��z:H��ށ���"#(e"�oE��ū��V��{��(���f11"t����H�)P� b*�?N��%I��:�^���U��c�j4c�(k
� �bt�h���Tc�F�
7���HWh�;'�/ѣ�N:�Ŗ���N�X~D����-�4g_�kD�h:5��g �+�Zt�6e2dȆδYFu���쓭F�vKZ!B��Ō�4*%i��l�e_	�����=�CBEV�B��,z=C����
B�	�h��!�Gz��+ ��X��W�.�ֶ���H���y��%��
�)��.���*�������Ë-ŪlbQ�c$����R� Җ��P���3�U�α���?T:��:u�,Z��R��,*@���k�EwI����FX� t��e�G�..k���k��֧X��4kZ2��B��#�� �Uk%��N:1о#d�L=]��V�����L���8@�����{�1��IU4s*�J�Z�,�#%by��Fө�	}���B�ۏ�����K�
� ��V��ȕو�H,h8�Fwz;�V��k	��9%�:q�'��;!�*��h�C�z7��Ю?q9�"
jeV2e~��q�t����-:LJ$����*%�e�C0�c�YZ����h�IS��d8얬X���$��+�	9*�r�X ��Y�T1%1x7�$��=����F�]@ Y�QO�XM]^ �@-���b�!@チp$���j����!"l=���� ��c��9����w�;�H��c�#G�aj� »���fb�ddى�B��u�ӭZuC��dֿNT��++�Es� %���3�K�e�f�����������J5��ş��8r���U]����-Z�4��:rј�����:�:�x	Qp ��Г��ÛRX��T���W}
9@_�CO�A��E�Kل����AE��wxs���u���Tf}��+�t'�,��)�T9d���{� �&�Ѵ:T�;���,���
8�����Z���w�!\N�0r5rR2��j���T���U��!��kaf(VY�cF�,���
��Oѣ~�b-4N�;%�ӭNt��_
�|N�����|��z"�w������b�b��Ĕ��cc�`	KS��j���k�r�+8ø��x�<�y� �jv;� �E�d"ƈ�cv;�׈����E� ,�\<$i�5��I_�
*Ŏ����S�ʡL��b�$�ҨZ!*U�ƋV�&M;�$�V�Ye���P������ǫ�U��\\\\\\\\\F�*��s\�_A�Wc������;$h֕:��¬�&Tq/�Q�?��n�"`H�F�PB6������z�IEB�	P����z^^�) ?&Z��LDDT�4(X\``(�`�O�%Hu9:Ы1
���� p*1R	ӲF̨�	ʽc�er�G�#F�c&�-GBM8�	�G�d��Bk��J*^��^��c'���W��W�B�u������τ��G *�
էSѳ-Gѣ��'Bt���Z4B%��J�a4�63�w�` d�	�F2�	x��,��m燆K�	�S`Ђ�V�0 �f��5 �4Rҗc��ѰZlj�,S)v���g �� `Cs̰9�,T�P��i�X�Wo{ul��L��\��֓WB�J�0�7�'J�f|:�:քɴ~������ѴhD*b�f�Z��`�?닋��������J�\���``w����U�/ΉX���J��1�[%�th]�V�T9W%p�� �z<Ao�G�(P������{2�R�"�� .�7�R&����QDC� ��
ll���Y6K��@�ADAĉT?&U�a$щ&�8���J��2~��>:vZ6H�=9ޜ���4 tu�ʩ�h�̟�q���z��H�UJ�	�$����ǥZ*V�~�G�oѣjՌ�~�v�P�:M� Ib�J������%y���BB�IKK^oV�J�%�<s^Q>UB͑q�A��c����v;�j��'bJ�Kk�1�� $��h�P�h+:+�hs�H��r��ZZ��w��)5;��
�����������g���]$֪T���VM	cfh�������G�N�Q�0�1$�����:�������R ^ �)�\Σ�<�Jo΂�Fz���k&M�z��d��#��)�Q�����$优#� <0��p���B� ��NC��KCN� b4^�*rAM�X Q�(��WX���qӝ*�~�uL��T4�c%B�h�&%!�tl��N�1�F�5�Q�F��,��ٙc����G�F����E��d�j5��,X�b��߿~���èd��:"tT�a/*��bz:rr��F�1�,d�:�C�Z��urS�Z�����K! �d�^��am����9c�e���l�K��]PR��B��M�k��@ @�,�K���/�p��8����U-�y�X��Enl�;�
�ȥ%/kȃ L櫬h�A�׀�[����R�*�(���b�l����d���1����>':A���ѣF�4k��4iв��FbJ�d���p�(�_\N���U�DM��ʛ�4)]A+M����p�o�Al��FAXߐTS&��%�k��%�FL���!\	�z��h���I5��@ w��	=:@1A�z�r
�~��Q ��La��R4��t��FU��B����ـ���,HN̮�~~��SW# ��%��#F8��Z�q֭ӭ��c�=�>��u��-B�k!*��TW~%�9Tl�2dɓ&HѣF�4mɝf*����M!^�$�w�HV	C��4hߎ�iQ"P�~�vIʓ&U;#���;�R#��-��R �	mE]y����T� ���c�!{"6��'��qz��������p� �8�*˧�N+��ԥ�< ��jj^oo]ul&���$�]�6�`s{e�
��)p������`���`V��&�*U;%�U��B�:թЉ|Wf*�4hѣF���F��V���i �D/���/2S�5qp��9��z�Y_���@eQjW�SrB@p9��C�Y�;�ӡ@�s��`�R�g�_��^�' ��mH�^ �WP��*Jm���%,"�7�9g��'G�����Sh�0��//x����+�*�L�)�R�f:$� őR��H}�F����#~�w�ߧN:4��B�6K�F�j��F�ѿ������{���Ы�~����߿�SH @���,4�9+w�#�[�h;�hѿbҢI�h�kE�Ήu:ŅH- �TU�$�(@h�e�
,4F2 �w�����;Yަ�.5�@F*�n�p��X0X�D�$�ѹ�4(`$Q��a������Sd���1A�ʪ�܊�.�(�4U-Rt������(z~@���.2.�*��2��&ƨ��	ӧN�hT�30�쑣F�4h�:4h�~;!�:�X��"uM��	c�.*������G��O�З�
,X��#B�B��; ���5r��:��y�W�].��h	��Q`i�#���9 }�i�����@� q(T�ɥ�,����G��������Aۍ$o4�Y$(4�i�2U��R�Gï�dtT=��zUP�~�1ΝZ�a7�gƈѣGߧ*�%���z?�~;D$ٖY2 $�!:�7���gZ,F9�E���'H�s�������h߲X�u��:%�	�$	:���eKΣ/
Zt��;�Haa`�(��� (<1x�(55�x�%��Mv5%�]��`dJ��L���8R̘�O���PWQ�W�E���G�e���T���88��y�����M��]ΐv4� l�b,z59�TAB�N��:TK⺻3�D"_�	�:$�����.thѭ��#�(<-!�n�(R�c�,r��?~�zR��h�ӝ/%Te��K���@!A�taa�j�Z!:�	��%��O��{B0�"] �i�$Ӆ��=W��K�*�l�C���
��d��Q��K��L_����5��	S/f:A�M��T|Tr��~�I�S�U~���Z�6GZ?up@D���N��qpw�߬ߣ:>���ӫ�ʪ�HfdUo��..W�F�\�"�hz��+q�F�qsG���Z���NtJ�I�u	4�gV��R�����<�.�ǈp�H���e�D�u,MAu)"9y���%%BDFzA���Yy�ɰ
�bE^M^,  VkAq002z;P���{;�|��x���9U��.��cS��t�����*F�6MVDWh�	4��Fc��':L�1'V�:T�E���.thѬ�0q�d���$��\\=*@�q��2#1QߴB�����G�x*-d����d��60B�f��h�����+�(�,�ad�O��P G�k���o]?H"z��,|}1���Z��(t�P5r�
� ��J��F,��FS�����=\�DT�LT��A�LN�d�1ߎʮM;&��#F�89�kGF���c2����6VL��i������&F$����.�������,�
���}N��>��������-N��E��~:��4h�i�ƈј��Z@�a�X�//w<�C���F�J Hs��� �	
#Hx;�T[Z�T��F�MN�
+�M�������y��dނ�4.�24RM,I$T\��U �Β�D	=#V fDv!��hAL�P��J� �����bt�ֲ���ѣG�֭Ό��C�h�\N�q9�L�b"��Ϊ*l�~te���>��H�c!α�T*ЪoНN�����ƜH����+�T`�QU<6#t�!�3�%2O�x�և/����T�N]&��`�	�jdG*d������zi��C2H�5�ʬ�j���u�� �f&��3�hН~��'닋�߿h�qqqqq�
�Q�X���'FA�K�3��v��Ϯ.�X�K�;"�rht#�,G�>�qߎ:ũ�!B�}t�ӧN�:��$�E��.!?9-u)?9l�W�^`�ȍ��s���,���R,w6^�g�n�R�W�b!���7�9�07=]����`eA��8Ul��/�גK��[��T؜MQ^ۏܣA
C $���J(�B�D^$-)ī��&��@�2d��2X�j�C��.th�я���o7��>�c�쉕\dM<r�����1/�硊I0�����d�p��X�Aѿ:ua21Zc�5�̱�PY��!�r^
�3]rM�rJ(c����)����tX�!�K�y��C�$�xl4b(�H
x�9�� �B�SW�DO�+� ����5�#t�ĭF�"jkѿG�.?F���f"/|*u=�q��ȟA��2ŶK��,\닋����J����О�\~��b�w�8�'h�kD�,Nt�ӧN�:�%{9���)����F B����|l�5EfWS&~�W%&��]j@ D)uEEz����V�g�k��0


�����������w��<JU�����%��CC'6�V$�+�#1�q��9)�-B$I�)�S�vKZ2X�jի�.th��#֧�fW: �4F���dwZ�|��6W�n��$�Z
r��9���ZY��4N��8�I��=h�u��)��fv��'<l��� �d�C�л�Q��)}%.�aGҡ�ldC��1�����(��D� �"�'0�3�Јaijih��,�/1w�+�*��^��t� tk�N���ӑ(ѓ"Xɒ�닚��������L� e�Bl���2����:θ������m\\B��* ����v255�ΣN��q��qr�tw�߿~��52qӲd���3���G�U	D�$:FA@_NTW������P$�&��-��2H	d$TI�V�J@"��p��k�b`�Ȼ�����l=���;�˓L�U�������A�/W�ev�V�� Qk�x����ru�ekʻ�rBu�_!X�0��F:�éΡ��G�X�	�����R�ҽYy(�Et���	e�"v���ʻڋ7쵍�?�B:�߿d90��G{�xJ��ps�՝U��w"����+������:NBƝ��hi��!�{�/P�x8ys���.])	"?##t����
��E�"���m
��D�T��(4vBTȀB��Xɢ���B�KP�\\닋���a���(^ G)��+H	���\h죤��
ɝ�g���d�գ�O�#d�w��d��ƅI�d�P���%�Γ&$�!$o���)�4bIFH���BC����"� Ȳ �Q(�P��J��<��  4�x�<ەR��)n���S�+Դ �� �|d�{RMM)`IVsP_/�-��`sdd49�Y��5���{@y�<^*�WQW���I�Z��jՌ�2d�a7�/��������1�B%P=��
uj����&c��8�� �5"�r��o��IBH����P����������t����#t���Lb�EDF�pY0�%1�p���� �`�00WhS�,�I���)� �x:@�]�*�!d�@�@
.�6�Q(C;p� xXX�D��D<Q��&%� ����5�ʳ$+�NɓB��u�����'ŕ��uE��G���.29"W �~r�:2e������Y\~����YGZ�:ŋU�#hD�t�7��N�dT��zz$�\� ��IaxPr����-����U]���l�;
Z�T���A��!�WT�Egp���J�����E)]g Mp��\+������
ή�D�6�V�s�F���4��
{Lkuy��;��@@d�to�߭h�:vH�:%�!����������hб�C�#3�л�e�(�t�������;\���gV�l��[�'�'!�1�gqt��h�hU:v53��X��e�z�aU!��ĥ��z�<�WI�(`xx��:փ���p@�A�AR'���1�(�V	"]u Pv����0=O��1�1�� 6�ށ�gP�:L��kS�N�:t�ߧ*Ҹ��,�Nu�:Տ��������'Y#x���������d�t9V��P�d�jՃ�X�:�K�:tJ��Q�P��!������E�A� �ߑ��"=^%�O����b�D�,�%s-9}6E���Q��	(���`E��A,VL`-E4`^Mx�����ÕIuYA�I� J�l���& �����UP)���}�v9�7��h�~:��"H>�d��=qqqs�?�k�B��0 �R�� l������`Y�,�x��ߕ&�n x�=^�Gcs�1�,M9�&�А�vc�3��d�P9�z"2�Vl���JA 
]� �!� ������b�Q��A��3�`\4(�T��(���@%111"
l�1&���< \��ُL@�!B � *A��'*lj�Qю�F����t��닋��k�}��h��7�Ѯ.?d�
rN��t���(��U�r��Y:ɑ�ʘ[0��V,�F��ɠ���d
� M ���!�� �H���D���FF�!CÅ��b�����DRl���.��Q���DC�[̝\!�� "T�ߐw������$���:�������;
E��Y�ٓUD_).�WT���<�0�ڐ���#e��&$��ѿ~;��H?#WZ���4u�����쑿:��B��!A͑��AAB �p��Q�����t��e`��N�8� `p��\a��, |tkD�1�������'ѣ��� 9�X�ZD.,*.Fb^2~�"1z=���T}������ADLB�_�@]ħ�ً�K��DO6��8!L�E��W#	t�K�H�v�D�ѿߎ:�"J���tk��ѣG��ߣ�d����4h�ӟ��*^"r^*J��z�1��D�cST1H �jŌ�:�;!։WWHW&$Jɫ��h���*"�H=*�c&�>p��Q\&�סc��5謚����{jv�6�S��
�K�P"$''#�l���+=^��J�k��%x�II�(�	x���6Z��OԊDFBQ�@����P��hY��!�K�֡$��V�N%]L�E��d;�u�����:��I�����w���� 3�W��\ E]@U ? 	w�:�Fb����c!�4&�~*̱c$c��G��L�D� �=�*D�|/HSc|z��:H�KBт+�������AI@_A�o�i�h������M����X�r2b��w*���F��8땨S� ���pttk���Q�F�\\B��z��k���k�������7�$"H�IOFC�J�?T|*����'�LT�!&��vK�N����c|Wf$�U�H$+�X�	׀(���r���S���)�j�{��[;e�r0Z�5_��[�.l�K���U�S�e�s8ak��T$Y�Z�nW��pj�ļ��� Īl\��ļX��g]`=Sy�����W�QU�Ƌ���@��X FJ�FtĈ�I'P�BTJq�!*�qӭX��?�?�=k-b�/�c# �b�`c��"$��..,\d���v�B���r�B:�����N����|/h����T��E^���&$�|c=1l����i��C�KӤ<DS��H#WW��Z2F@��
BqΣWN��ɋӤ�+�������������$�ɐ�A	�\\���$/��\\N:4k��οF�\d��2\��qqqq�$c�d����ߎ.��L$Qi苽��d\KF�G:���
�$ʴd:ӢD���2d��&�A�A$�*1�N�HX�YP�ȱ�kP�"�!��Գ����C��0�W�	k��( DD9�$�p�r�T�NWJ���Y���HsaU-5��s7N�D#3R��b��#ٓ{��R�y�QE�K\�(  ��Vvs�����4��v����+�om�������/B@Te�2dĝN�r	ߎ�vI�4Z�w����?F�gF�
�020Qg(K�+G�F��D���Ap]t�r:�������W2\F�A�MQ�H�����/#TAx�"��&X��x����� ^F*^rr�2z�ј�G�k��� ��K��H���F2
z��=H1W,H|����2���d���Ѯ#d�:�h�7���.......�ѣG��31�B�)+�SpҠC������2��2X^r�J̦"~�U�&KP�::��J�&Ls�
�:��$��߳=�:�]͗I2����р�H4	�� r�:���<]͇`�`ky`c�U�1�aѤ��Z04�4Zj��].<l6X��DAr�*�si��Ă��R�?X�p�:@�^�r��s$G��848D\你�m�+�U��M^p�=D2���B�A
�L��XT��&�u��-F��>�}m�!���4h���2X�hH�2��5�����������N�{p��\���L�]cK��A��, ƴ)� ؚX�h�r�}��@��l`d��].�0P��g�+���1��Fd��jd�'~��e^���9)�Cڐz��q�4:���c"kN�|:�#��ю�b��������h��4hѣ�Ρ�b�%9�z�V1�BW�PȊ�����*��� &�z�h:�bt�V�h���-
�B�aնDΉ 2�j1BR�F���p�"���]�KŮ�C����s��ف���.@ogA)@3y��� :���5=����J.�'���1M��D~*� nl�OY�QM����*�A�����%E���[.��w�x�P"B�y� ��^A�EJ��|&U��K�BL��d���-d�}���!���4h����kB� �3��#\\ �?\\w)�cv����g�"d�ƌQ�ht�ꨍ�9���uŝ��z�%l�]�/�o�U T��FO�]�l���_�ʕ:A��B1ı���Z���u9��Й1/�`mOd�gX�thߎ:?�������������������������4z4hѣF���M����B�Ɋ�����d�>>�u�ʜ���'*�u�-B�:ƈP�h�c"�Z-T%i[��ދ�!`�`/� �0��]؊��Z�"y��8E���E�n��M�
'ʨ�� dA`����� ���Xj����\���μ�JJ�	z��6X������j-0])s	,64p�& �`�J#R��J�������Pc��;� 	�Ujv�Y��N����P�N��T�iӕ&�q�~�t}r�4}�~�j�bk��qp�#��u;���eF��,'��j�F�DEoΕ�ƞ���=X�z��;�a����5 )x)���}
=X��"_ ���@�_�ɤ��H9S|T; D��C����U	�9Ve����N����th�닋����닋��������������4h��߿~�������T|Bz2 .F2D���m:'(@;�֒��@�F��h�b�$ӿ^C�h�r.�j �z
�Ɵ����8^�lJE�B�N� !��AQN[� V$!s�Đ=f ^�J�RPnujn3 y�9�7;݇�B��bk��yU|�kUVQQsM5ul��=�]�nV�!�#$�ơ��w���  j&�^x���6�G\d�`���d�aփ��	1���O��d:>�F�?~�~�`�ƈ���*���РǂC+�V�	?���N�TX��I�5�'&r�F�Nt���x�b���14��{�dI��������Td���x�4Z�"�}XU4i;2s�֫�F�a62hVZ?\dA\��#��:�����4hѣ߿~����ӧ*Mj1/�"t" ���}�B���i��XΒ��B��
��
�Z���P�h��%����us��A@�Њ�a�𔪠rj��K����`���2_5���×L̗�KUT\�Y�A��.�5u@w� CԵ5uU��,��X���ޚ�l((���^��TE䔕ӄ�$EdBR���
0Τf��iic!-�P�c`�(�a�!܊�Z��Ԥ�# Uj2δX�qΉ��e�F�
�Ń������4h�>��3�Dz���4oѮ.v22������ӧ~�C���~�*��r�x��
��F�_d̍hz7IjXb�x�a�R&I�6EU�4B;�H4\�X�Ҧ2��bJDJ�̜���U9�Gh������V2[�vKZ-��h�1��\\\\\\\\�ѣF�~����߿�g�&*�"�"͑�� z�EG��6��`��W�PqWŨS�Z��֋Z!:$�1"N������c#
w������<,h^���#Ol�hH&���*G��N�O˪�K��0b�{/y�����WW�\ڝI%�aY�x1����T�P^boV>KPv9A �	nV�Ų�6m]`v=^o	��tـXiX�01�TՀ�%��(��'I�*u��L�4 �u��e��Z=:��d:>�F�?~��d����(ߎ�a�yz͢�S̉���c*-Vg��P�,W1 ^* J���)��ID�;^c�����K��ȗ��4 �	ք�d�s?
9X,b~�th�2d~�,���qѮ!\qq��:���%����\\\\����4hѣG�F��4hѣF���@��p	R1��+��D%a��\f~����a��fF��
Ջ�BЁ���J�H%#|Z�iR0 ���-�	;2�k�#�Hs�Y�Z��j�p�hRA��k� �հll�.x��:����1����������Wcr�s:�keH�T��$1؊�|���4t&6[��P���W�s��L�&�� �6UPT�����O1F˄hhQ���2���*T�"S�f|Z����--d���w���G�(ѣG\�~��\z����3*)���IH� D] E���G�2��Щ��>�щ.R�x�:V^�`щʻB��֓1��ژ������*�Y��
�� 
2�T&$�:9���Q�U�b��..-GP�\��d����qqqqqqs������߿�F��4hѣG|#9WU d5����OZ���$s�n�q`�DrgV�hTH����6beP�ZT�Dędo��3�x�s�V��Š�����l�"�'F�fN�p�Ã�g�+����Z�x�:�$��<DE� /��W5P�c�ؘp�l�p��4�j\�.���P6l��9\̃m�A��F�L�%uP���5^{z$ "	u}��gy` �����A�%�
� A�E!	GƋQ�~�j$ξ������4h����W+������ߧx����fx�+����~�����M��u�� �N���W r�z;��@ �1r&L�wUA��J�:@��B�W-�LH��}:C�!�hQ���H�/���j�V?�Y!��M!Qnɕqqqqqqqqqqqqqqqqs��������:�mqq����x�VY'�%w��N�X��
p���]M��+��Q�fW{*u�r�N�*��li
�����ΝN�K�T(d��Oοx)��;�E�GGHf	sv);�F�Ň�˥�(�gH���@:��� ����T�����p����Ku&6Lo4	v:����U����˩H`9��Tw���T@J\�E�ГN�.29(����U���(Z���0���Q���F��9W�g��uG�)�ֳ���Z�b��ӎ��v��k�\\��F���_M)֫�~���������������qq'��o��B EN�?w��TЧ"c�����ܩ!/�7HK�2ըN��Y,F::ڠ �\$b6HLUʗ�#H����U��';32v6�������������������������eQ�������ѣ\\�*�+�T#=*�qq�����P�В��I� r�:�����8�	T-
�&$�Q$ĕ:t�5D�vH�d�;(`�ȗ�����ǀ(�B7�y(�80ٰ�y���i�,!�Wx��\�2 .2�l�^0�V20U2l��QBÑׅ�Ɔ��D0a��.�gM,x��� ����"�{�X���ըi��~�̂,�:��v%gW�B1�U�-��v6�����GdLH�d�[ZL��*��V�d�bգ��F:��d������?��?Z����r��~�qqqqqqqqqs��D����@Ñ�Y����,h �= &�1�f� �&�a�SP[F��o���M����BUa������Tur� �~DM����H1�X�v��GЧF�d�����������������s������e <q*��\\\G�C�v�닏�!f:b*M:Ҫ��J��� 'LC\-��AbS�B����VfHW �L���'V#�~�aց� /�N@@�'���G"z�6K[(�Lf��W���Q�,.�v:IW���dn��;z���.�jx  ���͖ ���u*��-]`l�"�����(F�FR֊hd,X�N:s��Ѫ>-x���Ce0�U$@��.���^o`a���a-O��P�:$��b_�4N%]jՌ�,Z��կ����\\c����h���qb����GF������������������������$bV���F��o  �W�`�a�B��]l��c��4/�H�GFu?Z@dDDd,�5��Ĝ���S#}����I֎U��qqqqqqqqqqqqqqqs�7��'h�����X>��t,�J渍��eOO_�ل�&%;�j�����W�$e� dN��xq��;���$�,h�
�J� ���L�1-	B��ևY�CIR^�L�#�E��3� ��I�������j�,Z��g{-Dv3��
[
@"��7Ap��ʂ4
��Z�R�I86_�j&fOmLFL櫭�s��U��EjJB�A����Phhy+���І���c9%*d�kl+:��6�(-ML��i�d�	S�S���htIխ�Z�jv�N�Z:ª�Y..����4h��;���!a�r��._�\\\\\\\\�\\\\\\�Ч�t�v�Ѵ?X�	��w��Wz	:�(��ZV-�X�LN�jӣ�T%?|B�� �~�?z�����XF"��������.�qqqqqqqqqqqqqqqsF��m��=�$e���W�������� ���QS�+D��Ty�X�̮F,�b-HN��E�_����B	ӧ:A��1$�!:��
sRmoT/ 2U`MuP5^g{M_ �T�Z����e"���f�U��mY���yʊ�@Ul);��륌�&��pQE@AIk4]g]`-K) :;'��0�1�t8<�U ,4U�!^Ek_�����"�IbH��TBbM����l�������C@�!&%�s��XU]�JçP�h���(S�*$�uA#������4h���qqp��ȋ�닗�.......���=s��P�hɓA(Y��,�X~FJ2"zѠ�d�td���I����@$�IP5D��{@1$O��ɱ��AFA�UK^��#�r�����(��1�����*���Qߕ9TN::x�h#xjc��uBl���B�FH��-&J�x�Cī�N����T�1'D��B��2P�NtJ�UOFKTڏ��]S'T����h4���u-Y�E��z8CF��T����\��E�/l���CC�יcp����J^`�˨�W7+� 	�h�0�-���l;%-CB"��`FA_\�����TC+����VG�C�-�JXpR�PPz&�OU�ي�dЫ$"J�*�FT�(P�*Uh쐡���M�e���?��~��qqqqq���?���#��8����wЈ�`�<ĂA�s����-�@o��4-:=�-���a�y+��D�^�.��������IH��މ�P'��5���Z�d����������������~�c����@4rB������6C�..�&r�^*J��~J�z*J�)W[Wf:�F�/B%:�
�|chU	�20����2bJ�d�jt�ʗ��^�f�'�h��V�T�FI�٬���A�̥%����0�g,l�9^�#MODG(h#���5I�p X�� {KH&�sz���\�םQņ��o��ss�H`!PP�(IhC���T�$ih�N�k�\!�.�o]v6�O�����a���	��ђr�Z���k�D�ӧh��գ�G�������?��..2Z:������7�����������R�ֿ�2G�HO֎�ƒh���4h��@$N⬞"�a�F,�S��X��*�b,�o���@k����̲�.�;C���"�hNFY�h�N�c�֭~�����������������u�G��w��G e�Rʐ#ZɡVZ֋��Ρ[M�.�x
��"��^����Y��O����x��TgV-BuP������(
�4-� �@K�T(J��K�ڒJ,CJȤE��
S畉x��a�����K��Eղ�j�d�����`dp4X�X,�*��\��0�x"Ʊ���7�9W�_a�[z[a؈�{oE_/3��6],�
_D�(] b��d�Á���iI��� r���`ˤ����h���P#8Y<�hS� Mm:Ռ�,Z����.�i��Z,Y���?���#\\\\*�qqqr�qqqqqqqs����~�q���6W������� ���,��Dr�Md-����o���l��&b�#x���@A@�N\�	ES�,x�FIB��d�]���􂬨�Zr�A:?���~�q��G�[�G�Lt*�w�Īl��'X�qqq
u���G�/��	�bj�R�Й{�ei7HdX�5�rDtuE�'*����@K�B�DbH+�*1�*M�Q��S�)�*넱$ؒ���	v"���5��
J�a4 9� ��p�ܤ�z���[۞��S��
����Z�X"�p�*������^�!�/6!��[{k	$�JUK�K�\.������.�EBWpPaK�u���rI�������V �b��P�Hz���F�{'I�`B�!�u�4#��U�q�ӕ:�`�kV4�������,NѣD㿮....-qqr������...................H�Ou���~�ߣF�4hѿ~�t����ѿ�~b^L�4�5r0S��@�d�^%�ŭ�xx���%B�r@E�:@k�����B4+Y��h?F9�����㿮#��?h
"&r.�8�c�5���$�g�IP CрW��`���X�x��/,l�@BF��N�d����w���'X��-
�|| L��2�#�*����n_�]]��@�����f��)l��FA�+�������#�Y4�5�u�x�Y|��9oEP/,l�Ş!"ȃN�F��BXs�a��q�+�����D9p��/p[��ɜ]�p�C�O��%�C1�3�"5%���XB��*DC	l莣 A�
���$ӧ&�@���H/Nэ!:4q��#*�����\\\\\F�������닋������������������bS���~�4hѣF�1ߣ~����i�'�Hhu ��GX�������d�:q'J�1x�>��""X��r
�	&����������������ѿq��?ӧ֬N�� ��_d����u�l�&LĔ�R�`{
x.�������F^�jz�J]]E�'B����t+H�v��ľ3BЫ�C�A����(�/�:�)$.�B^�K��&������gU-z��9E�L��US^����X��Jh)��A��\\ZR�/��+̰ ]�U�.��j%}Lŝʃ�%|w�ޮP��U� �j�r	��yi��Y��p�"��Ԛ�������jy�
<�댚!d�A�2$�
�	�����	߿닋��I�*u����F�F�qqqqq?��>���������������������uC�o��c���4hѣF;�o�NtH��6��#����ۅ٘ȟ�*8���@�X�@��N�^�*��I�(֏r���.#~8�\\\\\�e����z��ѿ~���c �Tq�u�tl��X��֋H���EQ���00`����� ���!�4�KA	fd�8���ɧd��662U�-d���5r '3Ueed%e�u��(#��u�D�A�ZH��4�՜Հ�������]�CeҖ�����D��z�4_"$�`�K�7���%�7���^ƕ,��BF��] ��RX�w�&��!`�B��q�q�Z�[��є�1�W��@h4��.Z�,�oU#9w��\�!��kGd���rS����j��!Ӵ�h�D(�q���3�����ߎɓ�����u���}qqqqqqqqqqqqqqqqqqqqp��T����ѣF�4c�F���������V=	3�D`Dq/������ѕŃ�B�)	A��E
���+�/t���\\\��d���������?�qqqqqsF���GZ�bƐ"��Xˬ[�Y U	�dʴcX�(2�gPdJ��t����1 ]22U~�����NL�ݑV3�i�>B�h�63�᭔�%��"�����.X�Ă���0UDv9�"���"�;�[Ɯ�y�/����y��� ���6R^
[�Rҗ�A,Mk<0Q�����M�$�EEW�#��Z�v�|е�@���,�.^�9z��78C��w�Ô�21�qK���L�,�4��Uw���!ѿh@���V�;D�h��Q�|X��5���w��֭X�jv�V�F�����>�����������������������fHfX�ю�4hѣF��4hѣ=z���كX�FY���a�dj�LH?�H�\\\p��:8
���l�jdaO�3l�4o��>����������������&C�=})���d��u��'X��!
�,ʇꄯV����Z�5��W/y�������7�����X�br�I�>N���H @��ߎ��A�7���;�a���X�Rx��7%��������59��  =����"�i_�ikRj�������RΠ��÷+"1*��A�j%��wV��@ '� �BI���h����ʺ|p����u<k8^R `z��/=��ԋ^��d�����h�
�p�[ %�i�����T|e��ET�'Z�+D)�S�Z�qq랍4kV�X�;D$Ь�5����}qqqqqqqqqqqqqqqqqqqqpvK����,�d�4hѣGF�>�aZÒ	ʌ))"�=<\(֔������*uh�H��XF*������ߞ��d@Y�̸����;��������Ύ����\\\������4h����ْ	R<�-��L���� bD�R]u-{ul�Ȕ�@�d��9[!��!��5vM�Z%]��Rdē|WHc|*��t�Z�~z�~��gM{z9@��� O_B��˩���+R�Bl����,.<fMrx7F�͗(`�c�(R����U�aA��S��gc�`�8�(dQl��=G �� �2V0<I4p��=�7�"8]
*�N�8S���u1�s� ���Qaz'`nl�L�ł���Zd.^b��z~��u��GI�:�j�ߡ:�bM	�Th�YF�vL�2w��d�9��~������...................#�B�9��#�F�4h��hѣ�~@Ix*��u�`�@ g�RV0��x���@�2���V5G�6a�E�ʝ z��(H��V�X�\G\\\\F�qqs\\\�F��t�I���=r���r�ʅ:BߣZ�b��c�T t��X8���:�
^�����y��Ō�cADd��_����-пdA �u5F2P�&~�t��꺡W��S�aAEy��v(<O�-1x6�E��W�T��O��["�]��}�J,MH&�oԵ��%g)��k�jcZ�+�qkd9Y�e�Aj[�Q�r#̱t(iUt1��dZ�x�p��-	M4R)2^z�8)��s�xp��iޤ,j�v�[Mؾt���]B^��/U �Ш�+$����3+�N����t��X�����G�#�F�w�ѣG�~;%��ߣ���닋��������������������\�I���G~�4hѣGѿ~��u5uB%21��VI��<%H>�����<�� �_�:ѣC��o�ǀ�C��A��y�닋�������������������������
���4F�]�����k�����\\d�ɒs��X;�2P󒮐��RU������
9� � �!�Ndo�H&L�1"J� U:ō	�	*�:t%D�����W=|

	1x;�
EILU����*:C�*�"<W�A��[Ze�`i���7M�@Mؒ��0���t��ʪ֚�,�ޠ`�bb�:��0���������6QW��D�e�l\���]o-)l�3�<RҦN*�����eqg+:�0Q�����PpVݦB��rW�a���j4�!)}�<_���t�3D$	�:v�βfS|h�q�,d:7�,d���4h�7�ߎ8�F��\\\\\\\\\\\\\\\\\\\\\\�q�\�R�N�~�q���o�F�k�6�V� ��r�%:�~;&c�22 'H`X�hK�OT�U��DIP�+�O&����7���N���3�v���-\\F�����ErT�$�ħX�iփ�d��D�]hxy*�F0�bC�4 ���(h�xr�P�b�``eQL�	�&$K1�|cUF�J�&�~ƅ�L�ѩ����*b��b�-	w
����A���]Α�����\|l��)VI_�u~��7��+$��(�6B���UG��Y*h�����2obI3U)Dp����L)ØJ�r��+9�₃r"[{��h��$�=����jg���H����w=���QT���AD@E�*Om�G5#�IAkԀꊇI�&�L�v7��َ�4WT&�`�X�to�,X����h��h߿~8�F��\\\\\\\\\\\\\\\\\\\\\\\F�q�\\d��e_�ɐ��ѣ�ߎ:1ΓBɕ�c�:�;C�p{�d��ru��B�x:�1Q,�f(�-\qju�Ѭe�\\\\\\\\\\\\\\\\\\\\\\\\�*�jύ*�q��P����_�j��X�'��@R�1SH*�iH���(*DD�"�j�"�|�X̱�����ɱ�%�PIT-!*%��kD��9uI
=SWЙ˥� �,s--uul 
�T�PL�^��Ii����G�	"��D��sz 01"��� B�QK�խ�%��r�9�$�K�P\���#I%,�D�&%�AaA��%d�T�A%�@]��QnRr�@��)��B��cW�aE��Vc��(*�{Ur��.��w;�ʎ�b�ʸ�eX���LU�X�ʱ���h�q�,d:7�,d���4h�4h߿q���G���......................_�;%��Ŭʌ�Y2X�c'�ߣ�o֣�Z:7����$`�H���p����	���