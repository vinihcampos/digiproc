3832
500
355
3
0 1
116 011111111
232 011111110111111
223 011111110111110
207 01111111011110
238 0111111101110111
241 0111111101110110
231 011111110111010
212 01111111011100
234 011111110110111
243 011111110110110
213 01111111011010
216 01111111011001
245 01111111011000
191 01111111010
165 0111111100
15 01111110
20 01111101
147 01111100111
196 011111001101
229 011111001100111
214 011111001100110
218 011111001100101
219 011111001100100
204 0111110011000
156 0111110010
122 011111000
18 01111011
52 011110101
143 01111010011
188 01111010010
160 0111101000
128 0111100111
182 0111100110
55 011110010
117 011110001
118 011110000
53 011101111
175 011101110
21 01110110
115 011101011
108 011101010
189 01110100111
187 01110100110
183 0111010010
56 011101000
22 01110011
23 01110010
174 011100011
101 011100010
114 011100001
57 011100000
184 01101111111
193 011011111101
205 01101111110011
247 011011111100101
209 011011111100100
210 011011111100011
239 0110111111000101
230 0110111111000100
222 011011111100001
217 011011111100000
63 0110111110
65 0110111101
104 0110111100
31 011011101
95 0110111001
136 01101110001
131 01101110000
98 0110110111
179 0110110110
70 0110110101
153 01101101001
133 01101101000
30 011011001
28 011011000
67 0110101111
173 0110101110
68 0110101101
178 0110101100
35 011010101
135 01101010011
152 01101010010
180 0110101000
29 011010011
172 0110100101
105 0110100100
6 01101000
1 01100
54 010111111
111 010111110
177 010111101
112 010111100
4 0101110
24 01011011
103 010110101
123 010110100
97 010110011
62 010110010
60 010110001
100 010110000
145 01010111111
197 010101111101
198 010101111100
192 01010111101
228 010101111001111
242 010101111001110
249 010101111001101
235 010101111001100
246 01010111100101
215 01010111100100
199 010101111000
110 010101110
121 010101101
109 010101100
5 0101010
59 010100111
94 010100110
99 010100101
61 010100100
130 0101000111
154 0101000110
107 010100010
27 01010000
26 01001111
25 01001110
176 010011011
64 010011010
32 01001100
8 0100101
113 010010011
58 010010010
102 010010001
106 010010000
13 01000111
45 010001101
119 010001100
3 0100010
2 010000
33 00111111
34 00111110
7 0011110
72 001110111
92 001110110
137 0011101011
132 0011101010
66 001110100
9 0011100
36 00110111
69 001101101
93 001101100
96 001101011
71 001101010
75 001101001
90 001101000
10 0011001
138 0011000111
134 0011000110
74 001100010
37 00110000
11 0010111
38 00101101
73 001011001
251 0010110001111111
252 00101100011111101
253 001011000111111001
254 0010110001111110001
255 0010110001111110000
233 001011000111110
220 00101100011110
236 001011000111011
240 001011000111010
250 001011000111001
237 001011000111000
202 001011000110
200 001011000101
208 0010110001001
225 00101100010001
227 00101100010000
185 0010110000
91 001010111
76 001010110
39 00101010
77 001010011
83 001010010
40 00101000
89 001001111
81 001001110
79 001001101
82 001001100
80 001001011
124 001001010
46 00100100
43 00100011
42 00100010
126 001000011
84 001000010
48 00100000
139 0001111111
140 0001111110
171 000111110
49 00011110
44 00011101
125 000111001
141 0001110001
149 0001110000
47 00011011
78 000110101
201 000110100111
248 00011010011011
211 00011010011010
221 00011010011001
244 00011010011000
194 00011010010
151 0001101000
12 0001100
168 000101111
186 0001011101
150 0001011100
195 00010110111
203 000101101101
206 0001011011001
224 00010110110001
226 00010110110000
144 0001011010
167 000101100
14 0001010
41 00010011
50 00010010
162 000100011
85 000100010
169 000100001
181 000100000
146 0000111111
148 0000111110
166 000011110
158 000011101
190 0000111001
142 0000111000
16 0000110
86 000010111
157 000010110
164 000010101
170 000010100
159 000010011
88 000010010
127 000010001
161 000010000
120 00000111
87 000001101
163 000001100
19 0000010
51 00000011
129 000000101
155 000000100
17 0000000
vinicius�U~O��}_���������^8���^4�4�ԍ��l�#e�)�E4�������������������������������hM)�E4���"�S@�hM)�E4���"�S@�hM)�E4���"�S@�hM)�E4���"�SB������%5�S_%4l���M|���M Cdl��j�v��(���x��1^;B�d#c#c#c#c#c#c#c#c ��� Cdl��!�6@��� Cdl��!�6@�h��C�v��!�;Tb�F+�b�F+�b�F+�b�F+�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b�b��ʡ�%�Q�%P�EP�r���-��m&�i4[I��M�h��E��-��m&�i4[I��M�h��Dh	F��h	F��h	F��h	F��h'Ƃ|h'Ƃ|h'Ƃ|h'Ƃ|h'Ƃ|h'Ƃ|h'Ƃ|h'Ƃ}�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#EF4 �Q�(Ƅb�b�b�b�b�F+�b�F+�b�F+�b�F;Tc�F6TceF6TceF6Tc�F;@����C�v��!�;Z�^Ԋ��v���F6TceF6Tce�nP|��&� "��E3ceF6Tc��rq�S|����rqFS*m&��A]��4�A>4�@Jԁ�5 jH.�h�4P	���	���	���	���	���	���	���	���	���	���	���	���	���	���	���	���pm�o�|����86���~"��{��86������z�_86�����pm�o�|������>	C��>	C��>	C��>	C��>	C��p'�|p'��C�C|p'�|p'�|p'�|p'��?��?�86����%�Q��	���	���	���	���	���	���	���	�p��p��p��p��p��p��p��p�p�
�p�
�p�
�p�Ѡ�Ѡ�Ѡ�Ѡ�Ѡ�Ѡ�Ѡ�Ѡ�jF�R6Z��ԍ��l�#e�-H�Q���Q���Q���Q���)�E4���"�S@�hM)�E4���"�S@�hM|��>M�&叓r�ɹc�ܱ�nX�7,|�w��|�w��|�w��|�w��|�w��|�w��|�w��|�w��6�#o6�#o6�#o6�#o6�#o6�#o6�#o6�#o6�o6�oW���'��>������������������
�
�jF�R6Z���[�M70#s70#s70#s70#s70#s70#s70#s70"�S@�hM)�E4���"�S@�hM)�E4���"�S@�hM)�E4���"�S@�hM)�E4��гr��r��r��r��M|��!�6_%5�S_%5�S@��� Cd&k\�,�v���pYL��W��z�W�F�>F�>F�>F�>F�>F�>F�>F��!�6@��� Cdl��!�6@��� Cdl��!�;@�h��C�v��!�;@�h��C�v���������(�v(�v(�v(�v(�v(�v(�v(�v5"}�6")�(�v(�v�˟#b&�O��E��-��m&�i4[I��M�h��E��-��m&�i4[I��M�h�"}��H�jD�R'ڑ>ԉ��O�#E�-H�jF�R4Z��ԍ�h���O���O���O���O�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h���I]�����Wci+�����J�m%v(ƄcB
1������������Q���Q���Q���Q���Q���Q���Q���Q��!�6@�h��C�v���v������1�� E3 �f��>M��r��ܠS0�`L���ܜ|����rq�5�7-�ظh+�\4F�|h'ƀ�h	Z�5�A�� ��=�ᡂᡂᡂᡂᡂᡂᡃ�>8�>8�>8�>8�>8�>8�>8�>8�>8�>8�>8�>8��J��J��J��J��^������(|�pm�a�^��J��J��J��J��J��J��J��J��J��>8�ᡂᡂᡃ�>8�>8�>8�>8�|����86��J8�>8�>8�>8�>8�>................"�.��^.��^.��^.�H�jF�R6Z��ԍ��l�#e�-H�jF�R6Z��ԍ��l�#e�-H�jF�R6Z��ԍ��l�#e�*1��*1��*1��*1�� E4���"�S@�hM)�E4���"�S@�hM)��r�ɹc�ܱ�nX�7,|��>M�&发����������F�m�F�m�F�m�F�m�F�m�F�m�F�m�F�m�f�m�f�m���W���'��C�>+��������-H�jF�iS1��0"�n`F�n`F�n`F�no�������f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�c\,k��p��5�ƸX��c\,k��p��5�ƸX���Z�Zf�f叒��)����)����)����)����)����)�ݠ ۴=5A3Zಙ !ڣ�1^��������6@��� Cdl��!�6@��� Cdl��!�;@�h��C�v��!�;@�h��C�v��!�;@�h��C�v��!ڣ�1^��1^��1^��1^4�B��г<.b�6�,�=3�@J�أأأأأأأأأأأأأأأ�ԉ��O�"}��H�jD�R'ڑ>�M�h��E��-��m&�i4[I��M�h��E��-��m&�i4[I���1^��1^��1^��1^��1^��1^��1^��1^�أأأأأأأأأأأأأأأ�; ; ; ; ; ;@�h��C�l��!�6@���)�E4���"�S@��� Cdl��!�;@�h�Q��(�d ��@Cb !��\�)�>Je�f�PY�TnU��O��s�\6">M��ɹ85�|�g���Ci6"
��h�#E�-H�m$�6�{HIR	"jD�����������������O���O���O���O���O���O���O���O���O���O���O���O��(|��(|��(|��(|�pl>	G|\40\40p'����a�J��J��J��J��>8�>8�>8�>8��J��>8�>...8�>8�>8�>8�>��J8�>8�ᡂᡂᡃ�>8�>8�>8�>8�ᡂᡂᡂᡂᡂᡂᡂᡃA]����W@h+�4�
�t������h;F��h;F��h;F���-H�jF�R6Z��ԍ��l�#e�)�IMjJkRSZ��Ԕ֤��%5�)�IMjJkRSZ��Ԕ֤��%5F6TceF6TceF6TceF6Tcd���"�S@�hM)�E5�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#]�5�#\,�`Yf��́e��6�l,�Y��R�%-�R�%-�R�%-�R�%-�R�%-�R�%-�R�%-�R�%,:��T��R��>����������������jF�R6Z���T�m*f6��n`F�n`F�n`F�n`F�����nXnXnXnXnXnXnXnXnXnXnXnXnXnXnXnX5�ƸX��c\,k��p��5�ƸX��c\,k��p��5�5�5�nXnX�)����)����)���nXnXnXnXnX;Tb���*1^;B�d�d#c#c#c#c#c#c#c#c%5�S_%5�S_%5�S_%5�S_%5�S_%5�S_%5�S_%5�S_%5�61�61�61�61�61�61�61�60v��!�;@�h��C�v��!�;@�h��C�v��!�;@�h��C�,�\nU(�vx���v[�Ae2����������������������������������h��E��-��m&�i4[I��M�h��E��-��m&�i4[I��M�����������������Q���Q���Q���Q���Q���Q���Q���Q������������������!� !� !� !� !� !� !� !��؉�61�6"|��|��|��|��|��|��|��|���M|���M|���M|�����&��77ɹ�M��S_%5�S_%5�S_%5�61�61�61�61�S.|�˟%2��L�,ܪ7*����魠&�<5�Mm�[@Y�TnU��O��PX�d,k2Y�|�g��ʦ�lDԎ���i+�����J�m%v(�v(ƄcB
1��O`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�O���O���O���O���O���h`�W@h+�.8�>8�>8�>8�>8�>8�>8�>8�>8�>8�>8�>..4�
�������������������������t��A]�vD................4�
�t��A]����W@h+�h;F��h;F��h;F��h;F���-H�jF�R6Z��ԍ��l�#e�)�IMjJkRSZ��Ԕ֤��%5��6���Ksm-ʹ�6���Ksm-����"�S@�hM)�E4���"�S@�hM)�E5�5�#]�5�#]�5�#]�5�#\,�`Yf��́e��6�l,�Y�,�`Yf��́e��6�l,�Y�:۠m���[t���� �n�uK|���K|���K|���K|���K|���K|���K|���K|���K�a�,:��T���������������ԍ��l�#e��6���KsQ�l|�w��|�w��|�w��|�w��|�w��|�w��|�w��|�w���c\,k��p��5�ƸX��c\,k��p��5�ƸX��c\,k��p��5�ƸX��c\,k��p��5�ƸX�,�zlzlzl	�0�s	�0�SC�hM��ۛ�kc�k`Af�Af�Af�:��
�!^S^�ZA� �nXnXnXnXnXnXnXnXSC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��60:l`t��鱁�c��M��;B�hX��c�,v��б�m�b}�+��#���ȯQ��cn���^��^��^��^��^��^��^��^��^��^��^��^��1^��1^��1^��1^;@�h��C�v��!ڣ�1^��1^��1^��1^;@�h��C�v��!�;@�h��C�v��!�����������)�������)����)����)����)����77ɹ�M��no������r�ɹc�ܱ�nX�7,|��>M��r��ܠ�7(��Ae3@u�<nO�iBf��3ZP��+г8�,��iBf��3ZP�rx:ܞ�'�Ƴ!cY���(Yf��5�(�e�H���Q���Q��!�; ; ; �J�m%v6��I]�����Wci+����ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԉ�jD�5"{�=�H�ƤOcR'���ԉ�jD�6�B
1]�WD�M5"{�=�ᡂᡂᡂᡂᡂᡂᡂᡃ�>8�>8�>8�>8�@J4�H�ƤOcR'���m&�I��OcR'���ԉ�jD�5"{�=�H��p�
�
�
�jGd���vA��p�p�p�p�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�jF�R6Z��ԍ��l�#e�-H�m*f6�3J���L�ҦciS1����T�m-ʹ�6���Ksm-ʹ�6���Ksm-ʹ�6���Ksm-ʹ�6���Ks)�E4���"�S@�hM|��>M�&叓r�ɹc�ܱ�nX�7,|�w�g|�w�g|�w�g|�w�g6�o6�o6�o6�o6�o6�o6�o6�o	�X0&�`M`����5�k�|���a|��a|��a|��a|��a|��a|��a|��a�a�,:��T��������������p؀�l@\6Z��ԍ��l��3KsQ�lQ�lQ�w��|�w��|�w��|�w��|�p�́e��6�l,�Y�,�`Yf��́՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��� ����Ǡ�Ǡ���s	�0�s��6�noA���6���DR�q����!� �rǠրAf�:��
�r��r��r��r��r��r��r��r��s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�r��r��r��r��r��r��r��r��SC�huM���4:��T�鱁�c��M��60:l`t����;B�hX��c�,v��ס�D4�Z���X���@^�7(��hX��c�,v��б�;B�hX��c�,v��б�;B�hX��c�,v��б�;Tb�F+�b�F+�b�F+�b�F+��h��C�v��!�;@�h��C�v��!�;_#c#c#c#c#c#c#c#c#c#c#c#c#c#c#c#c�d�d�d�d�d�d�d����ƸY�`X�7,�f�f�f�f�f�f�c\,k��p��Y�,�`Yf��́e��6�h�hVh��4A՚ ��uf�:�\Y���f��3ZP��+г8�,�=3���A�2m̄s/B��г8�,��iBf��3ZP���u�8m��g�#[B�ܠԍ���Q���Q����C�v��6��I]�����Wci+�����J�m%v5#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�#E�-H�jF�R4Z��ԍ�h�"{�=�H�ƤOcR'���ԉ�jD�5"{�=��Ђ�WD��6�BH�ƤO`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`�h`��"{�=�H���hA��m&�b�&�OcR'���ԉ�jD�5"{�=�H���������ƤvA��jGdI��h����h����h����h����W`�W`�W`�W`�W`�W`�W`�WcR; Ԏ�5#�H�R; Ԏ�5#�H�m*f6�3J���L�ҦciS1����T�m*f6�3J���L�ҦciS1����T�m-ʹ�6���Ksm-ʹ�6���KsQ�lQ�lQ�lQ�lQ�lQ�lQ�lQ�l|��>M�&叓r�ɹc�ܱ�nX�7,|��>M�&叓r�ɹc�ܱ�nX��e�ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ,��ͼ&�`M`����5�k�	�X0,⅜P��qB�(Y�8�g,⅜P��qB�(Y�8�g&�����XC�>+��p;E�d\6Z��ԍ��l�%5��6����k�ܱ�5�#\:�`ug��՜:��Vp��Yë8ug��՜:��Vp��Yë6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�8ug��՜:��Vp��Yë8ug��՜:��Vp��Y�444�[�[�[m�&�êhM��ۛ�k`��DR�)WV
��7�Hd �@:��h�tA6�+ރ[�[�[�[�[�[�[�[m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&�êhuM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SB�ki	Dk5M��Ͷp���j�HJ;B�hX��c�,v��б�;B�hX��c�,v��б�;B�hX��c�,v��б�;Tb�F+�b�F+�b�F+�b�F+�#c#c#c#c#c#c#c#c ��� Cdl��!�6B�������������������������������������������������6Vp�́՜:�`ug��Y�:�`uf��́՛�6Vl��Y�:۠m���[t�4A՚ ��uf�&ۮ	��m���n�&۪	��m�����u�8Y��˄�q�6�cХGz��B��R��
Tp�n0&ی	���2�ՙp�̸u�8m�[s���+�khQ��J��A�S@�����k䦾Jk䦾F�6�������m'ki;[I��N��v��������m'ki;[I��N��v��������m'ki;[I��N��v��������m'ki;[I��N��v���I]�����Wci+�����J�m%v�R4[I]�1��i+��#A>4�4�4�4�4�4�4�4�."�."�."�."�ԍ�h�#E����J�m%v(�dc�����Wci+�����J�m%v6��I]��.�A�4�A�ԍ��l�#dh;F��h;F��h;F��h;F��h;F��h;F��h;F��h;F���-H�jF�R6Z��ԍ��l�#eFnPQ�lQ�lQ�lQ�lQ�lQ�lQ�lm-ʹ�6���Ksm-ʹ�6���Ksm-ʹ�6���Ksm-ʹ�6���KsQ�lQ�lQ�lQ�lQ�lQ�lQ�lQ�l|��>M�&叓r�ɹc�ܱ�nX�7,�������,�Y�,��ͼ,��ͼ,��ͼ,�êXuK�a�,:��T��RêXuK�a�,:��T��Rއ��������(Y�8�g,⅜P��qB�(Y�8�g,⅜P��qB�(Y�8�g>+���p;E�d\6Z���T�jJkinm������7,|��>F��k�Vp��Yë8ug��՜:��Vp��Yë8ug��՜:��Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�8ug��՜:��Vp��Yë8ug��՜:��Vp��Yë8Af�Af�Af��kc�kc�k`M��ۘuM	�7�����n��\X*M��Af��h��|&���U���5�5��5��5��5��5��5��5��5�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�&��m�:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:lc�W��К� �� �����c�hX��c�,v��б�;B�hX��c�,v��б�;C��M��60:l`t��鱁�c �h��C�v��!�;_#c#c#c#c#c#c#c%4l��!�6@��� Cd,ܰ,ܰ,ܰ,ܰ,ܰ,ܰ,ܰ,ܰ,ܰ,k����p�r���nX5���ƸY�`X�7,�f�c\:��Vp��Yë8ug��՜:�`uf��́՛�6Vl��Y�&�DR�	�Q�u�6�pM�\m��u��@A`x �<X,��)��n0&ی	��m�ǡJ��)Q�A���J��)Qޅ*8M�m��q�ՙp�̸uf\:ۜ����W�f�kD�[�RS@��������&��)����)�1��*1��*1��*1��-��m'ki;[I��N��v��������m'ki;[I��N��v��������m'ki;[I��N��v����������Wci+�����J�m%v6��I]�A>ԍ�Wci+�����J�jF��O�vvvvvvvv���h����h����h����h�#E�-H�m%v6��I]�1��i+�����J�m%v6��I]�����v��x�W��x�v�h�v�#e�#A�4�A�4�A�4�A�4�H�jF�R6Z��ԍ��l�#e�-H�jF�R6Z��ԍ��l�#e�*1��1��1��1��1��1��1��1��������[�inm������[�inm������[�inm������[�inj1��1��1��1��1��1��1��1���r�ɹc�ܱ�nX�7,|��>M�&�cZcZcZcZcZcZcZe��6�xY���xY���xY���xuK�a�,:��T��RêXuK�a�,:��T��Rê[��c��c��c��c��c��c��c��`Y�8�g,⅜P��qB�(Y�8�g,⅜P��qB�(Y�8�g,⋆ȸl��ȸl����[�inj1��1��1��F���5* �@������M��o	��o	��o	��o	��"�m�7'�JǡJ��M��Ѓo6��o6��o6��o6��o6��o6��o6��o6��o)a, �����R�
[���k��D,iEO���azxA��xA��xA��xA��{г�;г�;г�;г�;г�;г�;г�;г�8A��xA��xA��xA��xM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘL�	��3\&k��p��5�f�L�	��3\&k��p��5�f�M��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`M�`uM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4&��m��5��5��5��5��Yރ[���5��Yރ[���5��Yރ[���5��Yރ[��,k�[xu��[xMK	�a6��)X�)X�)X�)Q=
TA����pAJ�F�h	�냫AՂ�ꕠ&�<X	���k�5)ǡ`e�X8��E�"����F�#X���k �5�a�3�ۊzqOCn)�m�=�����6➅*81"�X���3�5��Ĕ&�h��uK�`C]�na6� �n�����hM)�E4���"�STceF6TceF6TceF6TceF6@�hM)�E4���"�STceF6TceF6TceF6TceF6@�f�)�S0�`L�"��E3�^Ԋ��v���L�ɹ@,kD5�m'ki;[I��N��v��������jE{R+ڑ^Ԋ��W�"���H�m'ki;[I��N��v��������m'ki;[I��N��v��������Q���Q���Q���Q���)�E4���"�S@�hMQ���Q���Q���Q���������ХT�7,Q���)�cZ E4���"�S@�hM)�cZcZcZcZcZcZcZcZe��6�l,�Y�,�`Yf��͏�����e��6[t��6�pM�\m��u�6�pM�\m��u�՚ ��M�\�)U=
UA6�puf�:۠m��a�,:��T��RêXM`����5�k�	�X0&�`Ma	�!5�&�����XBkMa	�!5��q1�q1�q0 �@ �@:�`u"��E�ԋ�R,�XH��o=�'��D�7������"z�OCx�:�@:�@:�@:�@\6E�d\6F�3Ksm-�F5�F5�F5�F5�#\��#\ �T/uk�`m�&��m�&��m�&��m�&��&�m�B��6�m�B��6��70�o6��o6��o6��o6���5+jVԬ�X#R�F�`�a)a, �����R�
XAKzxAK
�P7�����E ���6��o6��o6��o6��o6��gzw�gzw�gzw�gzw�gzw�gzw�gzw�gzp�o6��o6��o6��o6�s	�0�s	�0�s	�0�s	�7��Ǡ�Ǡ�Ǡ�Ǡ�Ǡ�Ǡ�Ǡ�ǡgzw�gzw�gzw�gzw�gzw�gzw�gzw�gzp�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SC�huM���4:��T��SBm�&�ރ[�[�[���Yޅ��Yޅ��Yޅ��Yޅ� ��� ��� ��� ��
Xu��[xu��԰���,/B��B��B��B������pA`�F�T#X4B�PuJ�X	����W�`e�Xz^������A�\ �#H���(�7�1� � q 8�@�  � c� AJ�R���+�AJ�R���+��D��7�a���np,�<�,�(ƶ�i6_%�,��f��70�oz��Ƹ���M70"�n`E4���h���#s)�F�S@�hM)�E4���"�S@�j�l��ʌl��ʌl��ʌl���L�"��E3 �f�)�S0�b�l��ʌl��)�S1�nP|��I��N��v��������m'ki;[I��N��v��������m'ki;[I��N��v��������m'ki;[I��N��v��������m'ki;TceF6TceF6TceF6TceF6@�hM)�E4���"�S@�hM)�E4���"�S_���1"�&ۮ)�1��/�r���ɹc�ܱ�nX�7,|��>M�&叓r��� �� �� �� �� �� �� �� �́e��6�l,�Y�,�`Yf���|�w��,�Y�:۠m����u�6�pM�\m��u�6�pM�\m�=
UOB�PA`�#q��B�Sа\m��a�,:��T��RêXM`����5�k�	�X0&�c��c��c��c��c��c��c��c��`Ma	�/C��C��C�����5�5�5�5�5�5�5�5�Cx��o=�'��D�7������"z��iA4� ��PM"��)�IMjJkinm���ƶ(ƺ�k��Yf��͏��5���M���H�m�&��m�&��m�&��m�&��m�&��m�:��Vp�o	��o)a, �����R�
XAK�"5�F����#XDk�a)a, �����R�
XAK	��,�R0�FqB
XMg6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g�\ k�p��5��@��\ k�p��5��@�70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s70�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0�s	�0��5�f�L�	��3\&k��p��5ޅ��Y�� ��� ��
XAK)a, �����R�
XAK)a, �����R�kMKz�az�� �� ��p�ĨF�h��#���b�(�ĔF�J�,�/B��A�\ �.#H���(�4�8�"�#H���(�Ĉ`bD01"*� #H���/�4��"�#H���/�4��"��,ޅ��а{zoB���X=���`B�rǰ��Pu�8Y�|�k�c[�e��!e�ͽFno�sz�z��c\,k��p��5�ƸX��s|�����&��77ɹ�M��naf�f�f�f�f�f�f�f�Cdl��!�6@���/���)����)����)����)�f�f�f叒��)�Cdl���Q���Q���Q���Q���v��������m'ki;[I��N�!�6@��� Cdl��!�6@��� Cdl���Q���Q���Q���Q��"�S@�hM)�E4���"�S@�hM)�E4��Ђ��&ۮ�)�1�SBƴ�4O�r�ɹc�ܱ�nX�7,|��>M�&�՚ ��uf�:�DY���Vh��4A�� �n�u�@:۠m���[t��e��6�l,�m���[tjTA6�pM�\m��u�6�pM�\m��u��@��x�JZ�
�N)Dn#����M`����5�k�	�X0&�`M`����5�k�	�X1�q �8�zH=$�C��ă��A�q �8�zH=$	A�!�p�j�&�DH�	�Q�(�iA4� �EM"� �*7��⠃x� �*7��⠃x�:�h�Z��իCRS[Ksm-ʹ�5�����Q�uM|�p�R�%�Fno�s�B��B��B��B��B��B��B��B���6�Y�m�&�ë8M����#XDk�a�"5�F����#XDk�a�"5�F����#XDk�a�"5�F��� ���c�qDkAKzxUK
�aU,*��T���RªX1��x1��x1��x1��x1��x1��x1��x1��xUJ����U+�VT�
�XR�*�`1��x1��x1��x1��x�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�����3[f��l��#5�Fk`�����3[f��l��#5�Fk`A���A���A���A���A���A���A���A���M��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘM��ۘL�	��3\&k��p��5�f�г�;г�xA��x�J���, �����R�
XAK)b5�F����#XDk�a�/C��8�B�q0 �`�"��ĈF�DH�- ��E(U"��H�&B��T��D`�"�#H�����Q@Ĉ`�x�H�
�@V��P����=��PA����v-]��W`b���v-]��W`b�� �q8�@� A ��A���6⃦��cY����а2X�=�4�@�j�:��Vw�JǡJ�ɹ��p��5�ƸX��c\,k��p��5�ƸX��c\,k��p�r��r��r��r��r��r��r��M|���M|���M|���M|���M|���M|���M|���M|�К�Mf�:k@,ܱ�S@�ʌv��hM)�E4���"�S@�j�l��ʌl��ʌl��ʌl���䦾Jk䦾Jk䦾Jk䦾Jk䦾Jk䦾Jk䦾Jk䦾JhM)�E4���"�S@�hM)�E4���"�S@�k�ܱ�nX�7,|��>M�&叓r�ɹ`Xփ�ܰ���"��7,���u�cZcZcZcZcZcZcZcZ՚ ��uf�:�DY���Vh��4A�� �n�u�@:۠m���[t��e��6[t��5* ��MJ�&�D�)U=
UOB�SХT�)U=
UOB�SХTX4�G���ĊPbE(1"�F�<X4=�C��ă��A�q �8�zH=$�C��ă��A�q �8�zH=$	A� �EA"� �DH�$Q(��� �EA"�F�\#Z��W�OB�sе\�$Z���"��-W=	��j� �<o��⠂��A�TZ�-O=�ǡ�8�7����inm������1���e��65#dk��zH=u��[xMK�"5�F����#XDk�a�����6��j��Z�z{���Ū!�#XDk�a�"5�F���c����&L8�q0�`1���#XDk�a�"5�F�����R�
X�a�!, �����RªXUK
�aU,*��T�co6�co6�co6�co6�co6�co6�co6�co6�RªXUK
�aU,*��T����U+�VT�
�XR�*�`UJ�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6�co6��#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���p��5��@��\ k�p��5�f�L�	��3\&k��w�gzw�gzw�gzw�gzw�gzw�gzw�gzw�gzw�g6��o6���5+jV��#XDk�a�"5�F��Pc�qA�(1�8���0�F#H�#H�#H�Z�$W-�����8�$L��!�p��<�G7���W�x�Z�
�@?�����=�����H	�Z�7�����<�>��!cH�,o��"���9?�����-������-������-����1"�H��.`ċ�1"�H��.`ū�U��#X	���m�ǡ`\ �.H�	���"�Ep�z�ȍj��R� �@&���hu��[xu��[xu��[xu��[xu��[xu��[xu��[xu��Vp��5�ƸX��c\,k��p��5�ƸX��c\,k��p�r��r��r��r��r��r��r��r���Mf�:k@,ܱ�S@���Q���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|���M|��ɹ�M��no�s|�����&��70��5�ƸX��c\,k��p�́՛�6Vl��Y�:�`uf�ɹ�M��no�s�՛m�B�M�@&۠m�	���tm�6� �n�M�@&۠m�	���tm�6� �n�ХD�)Q=
TOB�ХD�)Q=
TOB�M�@&۠�)Q=
TOB�A`� �\X.,���� �h,���� �h	�랅*����F�<#q,�*��n��X.z����`��X.z����`� �Tq*8�J�%A���PAĨF�h�Zi�E�F�h�Zi�E� �Tq*�Zi�E��<Z�-O��S��P���Aj� �<Z�-O�Â6�(��8#o��Â6�(��8#o��m �H0F�m-ʹ�5�Q�u�,�Y�,�ciS_%��q H�8��,"4� Ū!�#XDk�a�"5�F����j��m�5�(�Ju%�/Co��k�a�"5�F����#XA�&L8�q0�`1��c���k�a�"5�F����#XDk�a�"5�F����#XB�XUK
�aU,*��T���RªXUK
�aU,*��T���RªXUK
�aU,*��T���RªXUK
�aU,*��T���RªVT�
�XR�*�`UJ����U+������������������������������������������������k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��5�F���q�#Y�����������������k8�g��5�F���q�#Yޅ��Yޅ��Yޅ��Yޅ��Y�� ��� ��� ��� ��� ��� ��� ��� ��� ��jVԬ,,,8�qA�(1�8���Pc�H©U#
�aT�*��R0�F#Z����T@Ū �x�*�TZ�
�O��!��ȱ�,o�B���^�?����y�i�@BƑ�X�;GazA�X�;�b��l^�-�R	��p� �!H'�D��H�i��"py�N4���8<�'?�����-������-������-������-��Ƙ� �q>���OB��Yfx�@B�үU���⠂��M��К�R�jXMK	�a5,&��԰�o���o���o���o���́՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��r��r��r��r��r��r��r��r�� � � �r��r��r��M|�гr��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r��r���5�ƸX��c\,k��p��5�ƸX��c\,k��p�́՛�6Vl��Y�:�`uf���5�Ƹuf��n�M�@&۠m�z���*'�J��R�z���*'�J��R�z���*'�J��R�z���*'�J��R�,������pA`� �\X.z���*'�J� �\X.���J�n%B7�����xF�<#q���G�n#�6�sХTX4�@A`��)U�u����PAĨ �Tq*8�J�%B4�@�"�#H��-4�@�"�#H��-4�@�"�#H��-4�@�"�#H��-4�@�"�#H����S�V�(U�Jo��Â6����8#o�Â6����8#oC Ɛ�1�2i�C Ɛ�1�2i��A�6�`��#i6���1���E� �6�xuK6���&԰��q0�Dq0�`1��c����&L8��-Q=�*�A6��p�
�Pz{��D�8���8���8���8���8���8���8���8���8���8���8���8��H��*��V��X_�<���+�⿎+�⿎+�⿎+��V��XB�Ua
�!U�*��T���RªXUK
�aU,*���?�?�?�?�?�?�?�?�ł���`���A�X �,x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��x1��T�
�XR�*�`UJ����U+�V�q�#Y�k8�g��5�F���q�#Y�k8�g��5�F��T�
�XR�*�`UJ����U+�VT���RªXUK
�aU,*��T���R�ŃŃŃ�$�$�y#$a�<���0�FH��y#$a�<���0�FH��������x�*�T�7��x��o�B�Ɛ���G������B�!i �@��X�;GazA�^�-�R	��p� �!H'R	��xQD�Q(J�S`|�l��zA�/H6��� ���`^�l����x�o���xy�O7����<<�'8����@<�s
�^���p���YJ�*�8,Q$�J���7 ���,/B��,/B��,/B��,/B�R�jXMK	�a5,&��԰��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́՛�6Vl���70��5�Ƹuf��́՛m�՛�6Vl��Y�:�`uf��́c\,k��p��5�ƸX��՛�6Vl��Y�:�`uf��́՛�6Vl��Y�:�`uf��́c\,k��p��5�ƸX��՛�6Vl��Y�:�`uf��́6� �n�M�@&۠m�	���tm�՛m�6��J��R�	��Vl���)Q=
TOB�ХD�)Q=
TOB�ХD�)Q=
TOB�ХD�)Q=
TOB�ХD#q"���H�n$B7!��ĈF�D�)XX X X #q"���H�������xF�<#q���G�n#�7���� �h��)A��7���� �h���G�n#�7�����xF�<#q���G�n#�7�����xF�<#q-O���S�ũ�b��1jx�<Z�-O���S�ũ�x�*�%C��HpF���m��xpF���m��xp*�.H
��R©�T�p�@�U \F����m �H)F5�c]F5�c\�`��T���8�$Q�(԰������q0�`1��c����&L8�q0*�@&�����C��x=����5�*�A�q_��q_��q_��q_��q_��q_��q_��q_��q_��q_��q_��q_�X�`y#P��X_�<���W��W��W��W��
�!U�*��V��XB�Ua
�aU,*��T���RªXUK?�?�Ńł���U+�XUJ���R�*��T�
�aU,*��T���RªXUK
�aU,*��T���RªXUK
�`��m���m���m���m���m���m���m���m���m���m���m���m���m���m���m���m�U+�VT�
�XR�*�`UJ����5�F���q�#Y�k8�g��5�F���q�#Y�k8�g��U+�VT�
�XR�*�`UJ����U,*��T���RªXUK
�aU,*���?�?��H�H�H�0�FH��y#$a�<���0�FH��y#$a�*��[��V�pUj��o��+��%7�C��{H�/i��#� B� ���#腤}���1{H�,Q'R	��pQD�/u'�J��QD�/Q(�M1��Һ�!GSd^�l�M�zA�/H6�Ƚ ���`<�'�����x�o���xy�O7����<B�O-\®'�c���=�� Ƒ�*��,��n�M�@�\H�=
V=
V=Хcа�а�а�԰��R�jXMK	�!,&��8ugzl��A��՝�5�:��h�xAf�M��h�xAf�M�@:�`uf��́՛�6Vl��Y���M��nac\:�`M�A�R�z���6Vl��Y�:�`uf��́՛ƸX��c\,k��p��5ë6Vw�������Yރ[�;�k`ugzl��A��՝�5�:���p��5�ƸX��c\,k�Vl��Y�:�`uf��́՛�6�xM���xM���xM���xM��
V=
V�xug�����pA`� �\X.,��B�ХD�)Q=
TOB�ХD�)Q=
TB7��P�ĨF�T#q*���J�n%A����pA`�F�T#q*��-4�@1"��JH�$R�)A��ĊPbE(1"��JZ��/�xd*�8H�$R��G�n#�7�����xF�<#q��)A��ĊPbE(1"��JH�$R�)BS�ĊP���1"� �<H�-O)BS�ĊQx�*�8i?��cHd�4�A�!�cHd�4�A�!�cHd*�.H
��R©�T�p�@�U�#i�AB6�P��m�F�RêXM`����5�kA�����&0�FqA�(1�8���Pc�qA�(1�8���Pc�qA�(Ua
�/��8��<���-XH��y#$a�<���0�FH��y#$a�<���0�FH��y#$a�<���0�F�8���8���8���8���8���8���8���8��,qE�(��8��X�Qc�,qE�(��8��X�Qc�,qE�(�`�c�,X0X�8�Ń�(�`�c�,X0X�8���8���8���8���8��,���b�#m�6�#m��*��T���RªXUK
�aU, k��?��pco8�$QT��R��XyK)a�,<����b��Ń�,,X0X�`�`�b��Ń�,,X0X�`�`��R��XyK)a�,<�����`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��R��XyK)a�,<����{�{�{�{�{�{�{�{�
Ղ�<�����#7��
� ��P�FH��-Q?�T@Ū �Hp<�4������z�P�D B� ҫ�Uc��D�!Q9�	���l(�-��E�{�<<�O���������aGSd^�i�M�z��u6E���QԘ/V6B���{�0B�?+�.��
��B�>��*��
��|�?
:����
��/H6����P4���lX�9֮b���X�{-_�Ĉ��j�q
��\G�#���bE�*�h
�V��n$A�����1"��`AK�"5�F����#qB��a6���m�,��
X1���co)`��R��� ��xA��;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;г�;���k;���k;���k;����� ��xAK6���m�-�Yކ��,�Cozw�gzw�g�X#R�Fۢ��m�!n�Fۢ�XR�
XAK)a, �����#XDk�a�"5�F�����)Xm�՜&���7���sХDX.,��k����<q8��G�n#�7�����xF�<#q���G�n#�7�����xF�<#q��'	�5���ȍjd�7����p�H0*�7����q�ȍjd �8H�$N'��ĉ�bD�1"p�8H����x]�o���w�.�7������
��i��A�i=�ǡĔ,�hzIBkT��ǡ�8o��­ �� ��$�Ă;��G��A�H#��w� ��$�Ă;��G��A�H#��w� ��4���H��4���H�mRêXM`����5��q0 �`A�����	A#8���Pc�qA�(1�8���Pc�qA�(1�8��<���0�FH��y#$a�<���0�FH��y#$a�<���0�FH��y#$a�<���0�FH��y#$a��q_��q_��q_��q_��q_��q_��q_��q_�X�Qc�,qE�(��8��X�Qc�,qE�(��8��X�Qc�,qE�(��8��X�Qc�,qE�(��8���q_��q_��q_��q_�*��V��XA�X1K��o
�aU,*��T���RªXUK������ ��m�Ċ!bEUK)a�,<�����R��XyK,,X0X�`�`�b��Ń�,,X0X�`�`�b��Ń�)a�,<�����R��XyK,,X0X�`�`�b��Ń��QR(�)B�!
E�"�B�D!Z�B��V�cy-a�<���+��R0�FH�ūŪ'�j�*�.
�UB���`��G����a
� � �Qi]NM+�l(�O
(��)�
A<B�O$Ŏ�����:��cL^�l�Ս�
��!W7E��ȽX�����{�0^�L����b��X�>+������B�>��*����|�?+��
��/H6����P������B�;���b��j�H�-_�Ĉ��"0*�8q
�R�G�����x*�<#q*,�n$@Ċ�b� ��#XDk�a�!W*�\P��m���m���m���m���m���m���m���m���m��m��m��m��m��m��m��m���,�B��,�B��,�B��,�B��,�B��,�B��,�B��,�B�#Y�k8�g��5�F���q�RªXUK
�aU,*��T���R�
XAK)a, ��xA��Ԭ�X#m��tB6���D#m�Ԭ)a, �����R�
XAK�"5�F����#XDk�a$W=
V-U��bE�F�TX.,�5�@1�x�<q8�'��ĉ�bD�1"p�8H�$N�IDn$�7Q�(�ĔF�J#q%���'kS"5����1�.o���V�c��J�8��$�C�+��J�8��$�C�(Ujd*�2Z�
�L�V�B�S!U����������x]�o���w�.�7����w� �#i��𸍤Q
+��pbA�G
��?������V+�B��!A���PyD(<�Q
(�?�w� ��$�Ă;��G��A�H#��#���??�#���?T��R�k����8��8�q0 �`A#$`��Pc�Z«XUk
�aU�*��V���Z«XUk
�aU�*��V���!H !H !H /i,o!�<���yk-a�<������Z��Xyk-a�<������Z��Xyk-a�<������Z��Xyk-a�<������Z��Xyk-a�<������Z��X��8��X�Qc�,qE�(�#�b�^���1zF/H����8��X�Qc�,qE�(��8��X�Qc�,qE�+�⿎+�⿎+�⿎+�⿎(y#$o��8��XB�Ua
�aU,*��T���RªXUK6�bE�"�����X�D,H�
�a�,<�����R��XyK)bŃ�,,X0X�`�`�b��Ń�,,X0X�`�`�b���,<�����R��XyK)o��8���8���8���8���8���8���8���8��X�Qc�,qE�(��8��+VV��X!Z�B�`�j�
Ղ��,o"��,o"��,o"ū�V?�V?�V�����s��*EO�x��7�E����^�/H� C���D�>V'����R��Ԡ>u6Φ��������ȽX����stB�n�ɁEq�Q\|W��Eq�Q\|V5B�ƨQX�
+��a��X`/VՆ�sT^�j��P���>_5B���\|>V�I�tB�n���
A<B�N��bƑ�^�>���Būر��-Q�Ū;��2�$L��S�T�P�E(U"�*�J#X4��ċ@1"��@ ��k�a�"5�*��V��qB�XUK
�aU,*��T���RªXUK
�aU,*��T���R�
XAK)a, �����R�
XAK)a, �����R�� ��� ��� ��� ��� ��� ��� ��� ��
XAK)a, �����R�k�a�"5�F����#XB
XAK)a, �����R�jVԬ�X#R�F�`�J�n�F�`�a�"5�F����#XDk�a�"5�F����#XDkUj��h��-�x�<�ġU����F�h��#�łP���U�p*�8H�$N'��ĉ�bD�1"p�8H�$N'��ĉ�bD�1"p�8#Z��L�֦A��pcx\*�
��� ǡĕ�q%$N'kS ��U�iV�B�S!U�����Ujd*�2Z�
�L��A��`y�i�A��`y�i��� �U`��01 �#i�p�x�Q
��?����� V=���a�c�yD(<�Q
(��B��!A���PyD(<�Q
(��B��!A���Py <�H$T��X0&�`MazLzLzL8�q0 ��0c�qA�(1�
�aU�*��V���Z«XUk
�aU�*��V���Z«XUkiU��Υ�E!
A{H����$o�F,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��Z��Xyk-a�<������Z��Xyk-a�<������,qE�(��8��X�Qc�/H���#�b�^���1zF,qE�(��8��X�Qc�,qE�(��8��X�Qc��8���8���8���8��,Z�X�`�j�bՁ�<���+�⿋?�?�?�?�?�?�?�?�֫��U�U,*��(��AU,X�`�`�b��Ń�,,X0X�`�`�b��Ń�,,X0X�`�`�b��Ń�,,X0X�`�`�b��Ń�,,X1�q_��q_��q_��q_��q_��q_��q_��q_�^���1zF/H���#�b�B�`�j�
Ղ�+VV��X!Z�^�0^�0^�0^�0^�0^�0B�"����"!cH�^�h���bA(� �X�2!H

(��* GS����ҫ�WS�\�[iU��*�=�V6Uca�V4��sd|�l��͐��0(�L/��������I�4��v�xnү�U�J�7iW��*���_4�� ���(�*
/���⠢��(�0
/U�J�0iW��*�ݮ_5ZUq�J�>+�����>u6�$�<B�N
4�b��B�;��A��y�,o���p�xd<��ũ�c���ĨF�TZ�
�OV
�jVL8�q_��q_��q_ŃŃŃŃŃŃŃŃŃŃŃŃŃŃŃŃk�a�"5�F����#XDk�a�"5�F����#XB� ��� ��� ��� ��� ��� ��� ��� ��
XAK)a, �����R�k�a�"5�F����#XDk�a�"5�F����#XA�������U�ł ł ��&L8�q0�`1��c����&L8�q0�`1`�Ujx�h��-�x�<�ġU��c��1�x�<H�
��\Gĉ��"d*�2Z�
�L�V�B�S!U�����Ujd*�2Z�
�L�V�B�S!U�����Ujd�7����p�H0*�
��Ă;��G7�­ �� �Q
:��*�E��Q|�i�A��`y�i�A��`y�i�A��`y�i�A��`U��,��w�� X�,W$�i(1 �H?�ă�1 �H?�Uac��X�~:�����c��X�~:������PyD(<�Q
(��B��!A���@0y <�H	�!5�&�����ǡ�����4�5�F��ֱ�Z«XUk
�aU�*��V���Z«XUk
�aU�*��V���Z«XUk
�m*�SJ�T>u.
(��F�yk1cy7�cy7�cy7�cy7�cy7�cy7�cy7�cy7�cy7�cy7�cy7�cy7���Z��Xyk-a�<������Z��Xyk-a�<����zF/H���#�b�^���1zF/H���#�b�^���1zF/H���#�b�^���1zF/H���#�b�^���0�FH��y#$a�<���1{x���@^� ,Z�X�`�j��FH���q_��q_��q_��qE�V�-"'��QbՂū���8��X�Qc�,qE�(�#�b�^���1zF/H���#�b�^���1zF/H����8��X�Qc�,qE�(y#$a�<���0�FH��y#$a�<���0�FH���k�b�B��V�
�!Z�+XQ�`Q�`Q�`Q�`Q�`Q�`Q�`Q�`��`��`� �� �Q �(�\!Q��TG�*#�E����DpB�!u����������V;4��f�\�ү��Ur{J�l5���\�iW�֕\��/�����\�?iW��E��&`>I��f+���p���֕�TҸJ�W	SJ�*i\%M+���I���16�&&>I���16�&&Ҥ��T��J�*i\%N4�S\�-k���*��|�j���P����W&4�ƛJ�i��M���<(�O����1z��^� ����qbA<�7�����H\*�8q
�R��S���UjxF�Dq"
�P
�P
�P
�P
�a�<���?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�L8�q0�`1��c����&L8�q0�`1��c����&��#XDk�a�"5�F����#XDk�a�"5�F����#XDk�a�"5�F��L8�q0�`1��c����&Pc�qA�(1��c����&R(R(\H��$AW ��UĈ*�DX X X X X X X X #q"���H�n$B7!��ĈF�DH��J��7��E+��8H�8�G���W������2�$L��!�w�.�7���������x]�o���p�H0<�4�� ��H0<�4�� ��H0*�
��� �� ��$��!A���H0*���S�XB� _=�����qbAX�G$ŉqbAX�G$ŉqbAX�G$ŉqbAX�G��H�H?TA��P ��X�/_>�W����� �:�TA�� �U`��0UD<�V+�������``�0yX�u??�������:���S���~O����u Oo���Q=����X^��	ikX�k�b5�F��V���Z«[��_���7�񼿍��o/�y���_���7�񼿍��o/�y��Ը(�DQ"���7�cy-b��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"�^���1zF/H���#�b�+VV��X!Z�B�`�j�
Ղ�^���1zF/H���#�b�^���1zF/H���#�a�<���0�FH��y#$b��{x���@X�`�j�bՁ�<���0�FH��y#$a�<�����%AD���F�8���bՁU�^���1zF/H���#�b�^���1zF/H���#�b�^���1zF/H���#�b�^���1zF/H���#�b�<���0�FH��y#$a�<���0�FH��y#$a�B��V�
�!Z�+X�k�b�(�0(�0(�0(�0(�0(�0(�0(�0^�0B�@B�@(�D>Q*i]MGRQ���Xp|�2ҫ���p��|�>V?���*���W>���f�\��_95����|��^6�sM�W4�U�u�^&8ׇ��Uܓj��f�+���p���ֹ�T�:ʜo�����q���o�7�M��q���n�7����#i\$M+���p�5�&��D�8H��	\�(w8J��L�Ɠ*k�f*��|�j���V�\��+�-r��ҫc�S`(�O
(����A�B�{��* �az�P� (B�/Q
4��ũ��xdX����!U���D�yj�<�To�����p�j�^� q q q q q q q q q q q q q q q q H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�q0�`1��c����&L8�q0�`1��c����&L8�q0�`1��c����&L8�q0�`1��c����&L8�H©U#
�aT�T�T�T�����D�$W?���Es��\�$W?��7!��ĈF�D#q"���H�n$@Ċ�bEp1"��\H�$W+���ċ@�Ĩ �\#q*
�R��S�T�Pc��U"�*�J�$L��!�p�Ըyj]�o��A��`y�i�A��`y�i�Ă8� �,H#��Ă8� �,H#�ZA��A�H#��p�PyD(<�Q
�L�����U��$�Ă8yD(<�/Q
���B��!B��z�P�D(^�/Q
���B��!B��z�P�D(<���'H��i]k`ă�е#i�ϭ+�l(�s
$��+�a
��B�v��E���z��X�,W +�����pb� �\ <�V+�������``�0yX�u:��@�ΠA5�&��	Б�1�#Z�kX1�`1�����o/�y���_ƒ�7�񼿍��o/�y���_���7�񼿍��o/�y���_��/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i/i,o"��,o"��,o"��,o"��,o"��,o"��,o"��,o"��!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�oo!Z�+X�k�b�^���1zF/H���#�b�^���DN7SC\�T!Z�^���+V�zF/H���#�b�^���1
Ղ�+VV��X!Z�B�`�j�
Ղ�+VV��X!Z�B�`�j�zF/H���#�b�^���1
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V��x��I
4��I
4��I
4��I
4��I
4��I
4��I
4��x�
AH�(�\>Q*
:����Uav�X]�Wk�����C�c�J�ҫ�5�綹\��/����6�|�ү����{�x�w$�mrM�ү��*���/��k��&`�p���eN�YS\�(q���o�7�M��"w<H��$�����������:����h�s��u�Z��\�k�#�s�u�p��β6��F�:��n�7����k�e4�S\�-k���*�ݮ_�����\�>W6B�ƘQ\�:����
��B�s���OaGS؅D B� !Q 
:���!BĂ8� �Q?B�������%Ɓcx�,o��@��T,iEO����D�-Q?�TO����D�-Q?�TO����D�-Q?�TO����D�-Q?�TAT�*��R0�FH©U#
�aT�*��R0�FH©U#
�aT�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T� ��&L8�q0�`1��c��T�*��R0�FH�H�H�H��$W?���Es��\�$W?���Es��\H�- ċ@1"�H�- ċ@1"�H�- ċ@1"�H�- ċ@1"�Z�$R��G����xd<���ĉ����Ujd*��-Q�Ū;��G7�����x(*�

����ࠫx(*�

������@0y <�H$��� ��g�~G��~$��� �b� U�o[�AV�PU�o[�AV�P�D X� ,Q (�@� �b� �D X� ,Q (�@� �b��m��D���l�@�QA��cH<�>I���kc��Qx�!_9�W�b�s��|�,W+�����B�p!b��\X�,W+�����B�p!b��\X�,V>����c�X�X^����H�kX�k�b5��A�%�o/�y���_ƒ�4�񼿍��o/�y���_���7�񼿍��o/�y���_���7���Zō�X�E�#�#))�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#��X�E��X�E��X�E��X�E��X�E��X�E��X�E��X�D+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�^���1zF/H���#�b�^���1zFҤ;���n��
Ղ�(� !Z�<���1zF/H���#�b�^��V��X!Z�B�`�j�
Ղ�+VV��X!Z�B�`�j�
Ղ�+V�1zF/H���#�b�^��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B�B�$(�B�$(�B�$(�B�$(�G��$>H0|�`� ��A��)-" �Ap�D�|�8ҫ����r�c\��WiU��U`�\��+���s�J�}/��U�sJ�Nk���5�aܓi��6�\�n����J�n�������q�K]β������q���o�7sĉ��"M��o4���x�Sojm�M�Q���"m�H��&����#�֍q�Ѯ7Z5��F��h�����������:�u��β�s��Ɠ*k���r�_5Z���\�?iUɃ�ct(�i��Ƙ�Ԡ!H'TNBS��X�Q
:���
�J�}
:��� ����0��(�~�B�ā�HdB�J!H%��R	D*#�����D�-Q?�TO����D�-Q?�TO����D�-Q?�TO����D�-Q?�TAT�T�*��R0�FH©U#
�aT�*��R0�FH©U#
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P
�P8�q0�`1��c����&L
�P
�aT�*��R(R(R(R(����UA媠��Pyj�<�TZ�-U- ċ@1"�H�- ċ@1"�H�V���S�U����Ujx*�<Z�
�O�B��xd*�8�7�E���8� �iV�B�S/���Z���Tp�x(<�
7���ࠫx(*�

����ࠫx(*�

���� ��`�@0y <�H$��Ƒ��i�� ��ab� �D X� ,Q ���{��X� ,Q $��Ƒ�X� ,Q (�@� �b� �D X� ,Q (�@� �b� �D &�Z�Ob�Qx�^9W�b�s��|�!_9�����c�y�<��(���رX�,W+�����B�p!b��\X�,W+�����B�p!b��\X�}+E���b�� ��ֱ�#Z��$�_��i�7�񼿍%�i"ƒ,i"ƒ,i!�<����BHC�y!$!�<����BHC�y!$"�^���zB/HE��!�"�^���zB/HE��!�"�(�@|�D!Q0<�_Ŭ<�E�$^���zB/HE��!�"�^��HHTL7��F�-a��,i"ƒ,i"ƒ,i"ƒ,i"ƒ,qE�(�#�c��R�|��^�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k4��D�"��H���@|� >i7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�
7�
4��I
4��I
4��I
4��I
4��I
4��I
4��I
4��I(�r��5rr��+�!i"��>QG�(�Ei]V��i]V�XƹԈB�@^�\!Q*
:��Í*���\1�_?5��r��|	ƾvk���5㛍|��_94�����@|�PiW���&�q�Si3�s���p�Z�U��-w:ʝ���M��"w?�Sok��M�	����0m� m�ě`q&�<�#��`�X�k�Mb0I�F	5��%��y��w<�o�m�x�;����"m�6�x&���5��q���n�6��P�p���3�&`Ҥχ�����1�_7ZU�d(�l���bp�\�V9U���P!{����>u>��O�GS�Q��!u?]O�P�z@`� 0^�,H��D-!�{xp^�����!�{Hx^�7���<�TZ�-U����UA媠��Pyj�<�ToEA��py�\o?�TO����DH��-Q?�TO����D�-Q?�TO����Dq"+�Ċ��"�<�TZ�-Uƀ��Pyj�<�TZ�-U����UA媠bEp1"��\H�$W+���Ċ�bEpUj��o�!��Hy�o�U@Ū �x�<�.7�������Pyj�<�TZ�-U��������D�y"x<�<H�
�R�R)B��T�P�E(U"�*�JH��ũ��jq�Z��ũ��jq�Z����x]�o��A��`� �,i��#�y�oG�cH�,o�@�� �� H $ � � � �@ y  <� �4��� � �@ �D�,Q=�Ob�P!b��X�{(�Ŋ'�b��X�{(�Ŋ'�{���^�/u���@��B�P!b��X�{(�Ŋ'�b��X�{(�Ŋ'�
��B�}�D*��
��B�}�D*��z��^�r����!z��^�r����!z��^�r����!z��^�r����az��^�v�����az��^�v�����az��^�v�����az��^�v�����a
��B�s���+�1�#Z�kX�k4�cI4�4����_ƒ�4�cI4�cI4��BHC�y!$!�<����BHC�y!$!�<���zB/HE��!�"�^���zB/HE��!�"�^����k�"*&�zBu ҫ�TL��!Q0B�`�D�
��*&TL��/HE��!�"ƒ,i"ƒ,i"ƒ,i"ƒ,i"ƒ,i"�B��V�
�>ik�K��Ƅڸ��k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X�k�b�B��V�
�!Z�+X��@|� >i4��D�"��H���`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`��`���HQ��HQ��HQ��HQ���$>H0|�`� ��A�����+�W �+Һ�D�B�G�(�Ei]V��i]V�XƹX��QD�^�\!Q*
:�Uq��\1�_?4���5�ۍ|	ƾvq���k�'��ƾrk���r�@|�PiW���&�q�Sn�s���p�8�f�7	k��T�p�8��n�m�M�Q���"m�H�F�Q�m`9l$�+@څhl$��6��m�8l�����k�p4�0I6�M����r0���M�F�o����z� M�	�jm�w?�\n�7��Ɠ*q�K\nֹ&`ү�����|~ү���sd(�l4����X�u-��BS��X�ҫ�Χ���|�}
(�OaGS؅��!H
��������@`��2!i�ZC"�ȅ �^�����!�cx�,o��@��h7���X�4Ɓcx�,o��@��h4���"��x�<�.��Ū'�j��Z���Ū'�j��Z���Ū'�"��H�+��@yj�<�<,o�T���X�J,o�T���X�J,o�T���*�TZ�
�UV���UAU����PUj�*�TZ�
�UV���UAU����PUj�<�To����UA媠��Pyj�<�T,o�T�ŪQb�(�j�X�J,Z�-N?�S������8�-N?�S������8�-N?�S������8�-N?�S������8�-N?��w�.i�A�Ă8� �,i��#�~4��Ƒ�X�?�@�� � �!H=�� � � �@ y  <� H $ � � �b��X�{(���B�P!{���^�/u���@��B�P!{���^�/u���@��B�P!b��X�{(�Ŋ'�b��X�{(�Ŋ'�
��B�}�D*��
��B�}�D*��z��^�r����!z��^�r����!
�lB�[���*�
�lB�[���*�z��^�v�����az��^�v�����a
��B�s���+�1
��B�s���+�1
��B�s���+�1y��y4�񼿍�<����BHE��!�"�^����BHC�y!$!�<����BHC�y!$!�<���zB/HE��!�"�^���zB/HE��!�"�^����Fo"������Mr�RmB�`�D�
��*&TL��!Q0|�D/H_ŬX�G��Mr�P�X�^���zB/HE��!�"�^���D�"F�F�F�*A\�\�u*
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�
7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�4��I4��I4��I4��IiRiRiRiRiRiRiRiR4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��I4��B>HG��!$#�|���+J���+J���+J���+J���V��k��q��k��k��(�D��uZWU�uZWU�V1�V1ƮA�W.:�TJ�����a����J�GiW��r��|	ܼsq��k�'r�=ܾOw/��k�Íx�k�m��M�ҸS�	�\�>q���n�ws����(q���������x�W����mz� M��&�Ǘ��&���+^�����>����>���+^M����+^M����+^M`:�6�_������n�p70I6�M��`�ɰq����z� M�F���G�����dms���u�4�ֹ&`ҤϚT���x�_7B����|�
+��*��
�l^�r���� ���(�r
+��Χ��Q��V����!B��
�^�/H��E�D�qHdB���E���{xp^���D-!�HdB���D-!�HdB�J/i�C���X�4ƀ��Pyj�<�TZ�-U����UA媠��Pyj�<�TH�$O�)E�T�ũ�b�(��2/o��T�ũ�b�(�jpX�J,Z�-R���W�J�7�_��+��%į�x��o��C��x�*�<H�-U���Ji�E��@�j�X�J,Z�-R��E�T�ŪQb��jpX�8,Z�-N��/�D�Ujd*�2Z�
�L�V�B�S!U���.�7���������x]�o���p�x(<�
7���#�~���� ���0��/i �@�� � �!iD-#� ��$_ă���}��A��H>��ЫH	�H>���� �Q;�N���yD�/Q;�N����D�/Q;�N����D�!u9�]NbS����!u9�]NbS����Q;�N���yD�Q;�N���yD�/V9ՎB�c��X�/V9ՎB�c��X�!W-�U�br؅\�!W-�U�br؅\�!W-�U�br؅\�!W-�U�br؅\�,W-��b�rر\�,W-��b�rر\�,W-��b�rر\�,W-��b�rر\�,W-��b�rر\�#o"6�i ƒ�7��H��BHC�y!�"�^���zB/HE�&L(�,Q0X�`�D�b����&L(�,Q0X�`�D�b���*&TL��!Q0B�`�D�
��*&TL��!Q0B�`�D�
���$B�`�X�|�D>V"+5��N��
��*&TL��!Q0B�`�Dƕ\�X�B����׍�Yƹ|�^���zB/HE��!�"�^���J����H�Q�`Q�`Q�`��@|� oooooooooooooooooooooooo>o>o>o>o>o>o>o>o>o>o>o>o>o>o>o>i#�>i#�>i#�>i#�>i-*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*A�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�+�Һ�r��r��r��r��r��r��+��+�+�+�W �W �W �/�4������|�8ҫ����v�xƼ{q��&�nI����x��_'�׊	��az�i��m7�1��Lk�g�s����j���鷉jm�Z�x���$I��5z�$k�mb0m�F5����Iz�k m����-�B�~ %<�������B��@�p��� Z8GX�t5�GCX�_�_���ޛV�Z�kլV�Z���Z$��5������z� M�F�o�s�u��q����YC��P�p���3���iRg���c\�LiW�����W'���r�J�N+�����m�u94��f�X�>V
:���E�QD�Q?TH�8�D�>Q#��C��D�p�@`��2!i�ZC!D���@�Q 0(�.H
$����ȅ �B�J/i�C���X�4Ɓcx�,o��@��h7���X�4�E�S�ũ�b�ོ2/o�ZB�����.!i�ZB�����.!i�ZB�����.o��C����y�8o��C����y�8,i��C�T�PbE��<Z�7�E�"��ོ8/o�Â��ོ8/o���"����.!i�ZB��`��!o����`y�i�A��`y�i�A��`y�i�A��`y�i�A�Ƒ�X�?G�z@0� ^�!Q ���@�� �� !H=�RaE �A�^�v(���'`��<�v(���'`��<�v��A�<�v(���'ac��X�s:��.�1��B�s���.�1��B�s���.�1��B�s���.�1��B�s��Ŏ�1c��X�s:�Ŏ�1c��X�s:��*�
�lB�[���*�
�lB�[���*�
�lB�[���*�
�lB�[�����8(�N
/������8(�N
/����b�lX�[+�Ŋ�b�lX�[+�����z�8^�N������z�8^�N������z�8^�N����$�A�$*����B,Q0X�`�!�"�^���Qz�/QE��D�b����&L(�,Q0X�`�D�b����&L(�,Q0X�`�D�
��*&TL��!Q0B�`�D�
��*&TL��!Q0B�`�X��W.q�Urࣩ
��GR*�pQԀQԀQԀQԀQԀQԀQԀQԃ\�T/HB����׍�Y��B�`�!�"�^���zB/HE��X��u"iTH�
4��I
4��A�F�i!F�i!F�i!F�i!F�i!F�i!F�i!F�i!F�i!F�i!F�i!F�i#�>i#�>i#�>i#�>i#�>i#�>i#�>i#�>i#�>HG��!$#�|����EiTV�EiTV�EiTV�EiTWB�H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ���EiTV�EiTV�EiTV�EiTV��k�V��k�V��k�V��k�V�ԉ�u"k�H��R&�ԉƬ\�W*M���R&�ԉƬ\�V.q�;�ʝ��Mr�S\�<ҫ����.5�ƹx)Ɠ �I�w/Sn��M96�P^��ԛMz�n��4��M1��>q�ڮ7[U��7M�KW��s�M6�"^�Z�tj�6��6��M�8�P�z�
׫l�w�E�P�_�	O'�r�y�.�Hr�t�*wHr�t�*wHr�t�+Hr�t�+Hr�t�+N�RM@�$�RM�)����)��-����>�b���+^��h�ly�F/^׈�m�M�Q����&��5β���`�8Z�s���I���mֹ&�iW����@|�Pk��r�A�W'����|�>_9���6�|�>V+4��C�Pa�0QD�Q?O�E�Q�((�~���)B8��G�O�GP����(�Q?B��'ࣨPQ \(�.H��D-!�Hd^���-!�HdB���D-!�HdB���E��zԸ��!o[��F�(�#�Dp�H�i"8Q�G
4��F�(�#�Dq{H�/H�����{H�/H�����{H�,i�������Ըy�2,o�-!qH\B����-!qH\B����"8Q�G
4��F�(�?��x�/i��#�~4��Ƒ�X�?G�cH�,i�� ��az@0� ^�/H���Ƒ�<�H$Ob�رD�/u(�Ŋ'�bA�^�v����'a��B�s(���'`��<�v(���'`��<�v(���'`��X�s:����!z��^�r
+��� ���(�r
+��� ���(�r
+��� ���(�r
+��� ���(�r���*�
�lB�[���*�
�lB�[
/������8(�N
/������8(�N
+���<(�O
+���<(�O/�����@|�P/�����@|�P������z�8^�N������z�8^�N��+��
�<B�O��+��
�<B�O������z�8^�N4�cI
�!T�<��L(�,Q0B��TQ
�!QD.�����TX�L(�,Q0X�`�D�b����&L(�,Q0X�`�D�b���*&TL��!Q0B�`�D�
��*&TL��!Q0B�`�D�
��Ur�|�Ƽhk�ʂ����D��� �� �� �� �� �� �� �� ���\�B�`�����\�ƼhiU˄*&TL��!Q0B�`�D�
��*&8Ջ��R&�D�Q��HQ���$>H0|�`� ��A����$>H0|�`� ��A����$>H0|�`� ��A����$ҤҤҤҤҤҤҤҤҤҤҤҤҤҤҤҤҨ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*�Ҩ�*��H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ��B�H\i�!q�.4�Ɛ��BҨ�*�Ҩ�*�Ҩ�*�Ҩ�*��:�s��:�s��:�s��:�s��V.k�H��R&�ԉ�u"w+�/W��ĚW�s�X�Ƭ\�W*w+�&��	��C�|yƮJ�/��׃��N4�s��6�v^�\׮��=z�l5��X�Lm�'��z�?^�����t���z�-^�
��aB�F�F���F�ZH�+G�������>�2�~�-�S�@Jy<×C�Cp7��I��RE�EHXT��β^u��������;|.�������o����R<���X��������@Jy	O&�h�m�����> �`q&�I�x5����z�$M�Q����P��;��7Y����k�'�7
c\�n��6�\�i�׍���/���\�OiW��5�|�ҫ�Us�\�}iU��U`�X |�>u:��A�Π�E�QD�Q?R�)AE�QD�Q?O�E�QD�Q?O��8�D0|�>Q
$����Q \(�.H
$��D�p�@`��i"8Q�G$���C䀡�@P� (|�>H
$���C䀠���(�~
(���'ࢉ�(�~
(���'�{H�!H

(��Π��P`���B�/i�D���@`Q 0(�#�Dp�H�i��C䀡�H|�4��� a�HB�!H���� ��az@0� ^�!Q ��T@* 
� �D B� H$@� �P!{���^�/u���N������!u9�]NaEc����,u9�Nb�S����,u9�Nb�S����,u9�Nb�c��X�/V9U�br�QX�V9�AEc�QX�V9�AEc��\�>W-���c�r��\�>W-���c�r�Q|�_'��E�pQ|�_'��E�pQ|�_'��E�pQ|�_'��E�p�|�>_(�����|�>_(����J�l4���J�l4���J�l4���J�l4����x�!^'�W���x�x�!^'�W���xQ&�I�jD��Q&�I�jD���|�/_'�����p1��Hy!$"��&Qc�!QD*(����TBꏝQ�/VE�ȽY�"�d^��Ցz�/VE�ȽY�"�d^��Ցz�uB��Q�
:�GT(�P��uB��Q�
:�GT(�P��!QB��J�@|�`Q���GU�W uB��Q�
:�GT(�P��>V0|�`Q�
:�GTB��TQ
�!QD*(�E��B��TQ
�Ҩ�iTH�
4��I$Ҩ�k�H���$>H0|�`� ��A����$>H0|�`� ��A����$>H0|�`� ��A��T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�U�QZU�QZU�QZU�QZU�QZU�QZU�QZU�Q]�+�Ew(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��QZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�u\j��r�s\�\Ҥ5�%ɵq�xq�p�w+�Ƈr��ܬhM��&�Ǘ����Wr��x1�^
q�ߝ��۬���p�����֠�8Zm����8O�g	�X�j����X�0M�L�ֱT�^�����`:5�|	5�&�Z |=^e���%<�"Sɿ�]�� !�5;�X�O:���VM�
�,v���� *h��� *h��� *h�y΅�4�SO3��<�U��Y:O:��yԎ�Τy�+�r�j.�)��-�B�~�>�c��|����<�#�������6�#M���7ĵ��-w?��n��\�?k�g�+�1��Lw$�n�MƼl8׍�MA�^'�������\�sk��mr�٥W>��綕X�V iU�U`�X�V :��A�Π�E�QD�Q?O�E�QD�Q?O�E�QD�Һ�4��M+�P�D�>Q#��H�D���@`�D�>Q#��H��8�D�>Q#��H��8Q�G
7���0��>i4� *@J� Ҥ 4� *@J� Ҥ 4� *@J� >u
+�����E``��0QX(�i�B�U�۹���p�4��z�P��>H
$���C�0��>i�@�*@J� Ҵ�m+H�Ҵ�m+H�Ҵ�aD��Q �!H=�Rb�؅ �!H=�Rb��QD(�Q
(�@�� AE ���D X� ,Q=��@��B�P!
��B�}����'a��B�s��� ��l(�[���{�l^�[���{�l^�[(���'!{�l^�[��*��
�8B�N+�����8|�N+�����8|�NiU��*�=�W'�����\�ҫ��Ur{J�O/�����@|�P/�����@|�P/�����@|�P/�����@|�PiW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�
$�D�`(�lm��M�I��6�Q&�
$�D�`(�lm��M�I��6�Q&���+��
�<B�O4���HC�(�D�c�,uE�ȅE��TB�]Q�>uGΨQ��"�d^��Ցz�/VE�ȽY�"�d^��Ցz�/VE��Q�
:�GT(�P��uB��Q�
:�GT(�P��uB�����H�E
:�GT(���N䚠��uB��Q�
:�GT(�P��ҫ�w/���
$!��!i"�|��TQ�!QG�(�E(��|���P�I
$#�WU�u"q��$>QG��Q�A��|�`� ��A����$>H0|�`� ��A����$>H0|�`� ƕ ƕEiRiTV� ƕEiRiTV� ƕEiRiTV� ƕEiRiTV�EiTV�EiTV�EiTV�EiTV�EiTV�EiTV�EiTV�EiTWr��Q]�+�Ew(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��u]�+��w(��Uܢ��Wr��u]�+��w(��Uܢ��Ws��+.�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�u]��N5b� ��H"k�K�j�ͲLȁ�1ܬhw+��ɵrTڹ+�|qz�8�_q�8���r�3�&��{^�ݗ�5�9�u�5��l�n�]m֡�|�:Ϛ�[U6�j�^�ׁkX�*k��q6�u�V�5��F��$ Z�W�h�t�O'�r�o�C�Cpn�"�y�+I�R7�*ȰQ���Go���Tv�]Q��uGo[��ދ�V����x�k���׷��t��GH
�t��������o����:O:�@CS��C�JI	O&�h�m�����m��V��k��ׁX� ^�	o4�����(q�KSo�s����j�γ���~�p�5�6�&�w/�5�aƼl8�j��{�|��W'5��6�\��/���s�\�{k�ϭ*�\�}k��m*�J� >u:��A�Π�E�QD�Q?O�E�QD�Q?O�s�3\�~iTO�+�SJ�~(���C�8� (|�G$�H�䀡�|�>H
4��� a�H�H iR T��D��(��T�� �H iR T�� �H 
(��OaE``���(�u=��������3��G���k�6���?��i7�
� yj\(� Ҩ��T�� �H iR T�� �H iR V��i�V��i�V��(�{��)�
A�B�{��)�
A�B�{
(�@�� AE ��QD(�Q(�Ŋ'�{���^�!V>�U��c�D�!u9�]NbS�QX�V9Kc�bp�Զ/u-��Kb�RؽԶ/u-��Kb�RؽԶ/u-��Kbbp�X�!V'��Erx�X�>V'����bp�X�>V'����bsJ�OiU��*�=�W'�����\�ҫ�����@|�P/�����@|�P/�����@|�P/�����@|�P/����x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���M�I��6�Q&�
$�D�`(�lm��M�I��6�Q&�
$�D�`(�lm�
�<B�O��+��c�,uE����:��TB�]P��VB��QYiU��YiU��Y
+!Ed(�����VB��QY
+!Ed(�����VB��QYiU��YiU��YiU��YiU��YiU��YiU��YiU��YiU��Y^����sy����%�^ �#4���H�]+��t|�����>WG��J����\괪�\괪�\괪�\괪�\괪�\괪�\�Ϋ�\�r��5cj�\�Ϋ\�ΫJ���+J���+J���+J���+\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ�Ew(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��Q]�+�Ew(��6�b�X�l�\ I�<�ɷSn�&�LM���u16�bm��۩��e6��Քں�VSj�mYM���e6��Քں�VSj�mYM���u6����m]M���u6������V\j�8Ռw+�w+�M��&�Ȝj��5r�r�r�S�\�6�hq��8�ǝ�������bm|16��I��W����Kԛ۹���I�M�_W��f���u�5���=��l&�-�s���:Ϛǁ�X�7^�Z�aSX�(m��ڀq֡�H Z	C�����m��V�h�y�.�Hr�y�+�"�t�u#�� *h���3p:�S^�CZ�ck�1�N��6���6���6��hm]1�jN�S�:�B��jo�9��������] +Z�N�3�޷��z�VN�
�t�V�]y���"�,*v�JI:KG�Jy�)��-�����5��b0m�F��ֱ�D�<�����Z���_��[U6�j��g��	�m&��^7\k�Íx�k�����{�|��_'���N5�x��+����\��_;8��mr���W>���֕X	�V:��) ����3\�{k��aE�>u:��Oc�Pa��|�>u=��A�Χ��0���>u:��Π��S����>u=��Oc�S����>u=��Oc�S����Q 
(�@Χ���|�{iU��U`&�X	�Vi]O�*�J�}iU��WS�J�Һ�ZU`&���ҫ4��֕X	�u>���M+���Vi]O�+���u>���֕��Һ�G� C�!��D|�>Q(��@�������(�Q
(�@�� AE �A�(�v
$��'1�ͥu94��&���V9ՎB�c��X�/V9ՎB�c��X�/V9ՎB�c��X�/V9ՎB�c��X�/u-��Kb�RؽԶ/u-��Kb�RؽԶ>_(�����|�>_(�����|�W'���ErxQ\�W'���ErxQ\�>_(�����|�>_(�����|�W6+昅|���aE�d(�l�����ҸSW
cJ�Li\)�+�1�p�4�ƕ�p�8�)�7
c��p�8�)�7
c��x����7e�I�������<|�O/��M�I���M�^6U�`|�P/����x�iW���x�iW���x�iW���x�iW��
�<B�O��+��c�,uE����:��TB�]P��VB��QYiU��YiU��Y
+!Ed(�����VB��QY
+!Ed(�����VB��QYiU��YiU��YiU��YiU��YiU��YiU��YiU��YiU��Y,	B�;���<���ۭSJ�`Uk4��>WG���]+��t|���ֹ�k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�Wr���sjˍYk�V��k�V��iTV�EiTV�EiTV�EiTV�Ek�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��k�V��w(��ܢ��Wr��Q]�+�Ew(��ܢ��Wr��Q]�+�EM���u1ܢ��L^�m�˚�⧙�y6�bm��۩��Sn�&�LM���VW���}^����z��W����_W���}^����z��W����_[e��_[e��_W���}^����Ƭ�՗���r�b�ڹRm\�6�T�_"w/�;�ȝ��I��Bm|��_w/�׆Skት�:�x)ܼ�^
M� &׀�0N�$�M�z�sknMc�9�u�5�������So������F5 孲���(m���`q6�t@�F���Ѐ@�y�OV���j	N�)��]0Eb�<�F�Y7�*Ȱ����t���􎦽�6�����N���Ö�Y[�eӵ3�jf'N��N����;S1:v�bt͠��Ae�6�Ⱥu���ږ
9��(�h�kސ�zJ;z逩�u�o��İ���)$��I'���-B�~�>�B����6��b0m�x��ֱ�D�x������Z���_��[U6�j�\'ɴ��m&��^7\k�Íx�M���{�|��_'���N5�|��+����'r��Ʈsq����s�\�}k�ϭr���ViU��U`�X�V iU�U`�X�ViU��U`&�X	�ViU��U`&�X|�{:��Χ���|�{:��Χ���|�{:��Χ���|�{:��Χ���(� Q :��Χ���ViU��U`&���Һ�ZWS�J�}i]O�+���u>���֕��Һ�ZWS�J�}i]O�+���u>���֕��Һ�ZWS�J�}i]O�+���u>���֕��Һ�ZWS�J�}i]O�+���u>������X|�}:�GΧ���|�}:�B�`�A�|�s(��WS�J�ri]KaGR�QX�/V9ՎB�c��X�/V9ՎB�c��\�!W-�U�br؅\�!W-�U�br؅X�!V'U��bp�X�!V'U��bp�|�>_(�����|�>_(�����|�>_(�����|�>_(�����|�>_(�����|�>_(����|���b�L(�l�����>I�G�6�J�Li\)�+�1�p�4�ƕҸSW
c��p�8�)�7
c��p�8�)�7
b��~��8�-��&�iRj��x�x�Ҥ��M�I���M�I��U�a�^6����A�^6U�a�^6U�a�^6U�a�^6U�`(�P
$��5 �M@X�Qc�,uE������T(�����VZUe�VZUe�VG���]+��t|�����>WG���]+��t|�����>WZ�u�WZ�u�WZ�u�WZ�u�WZ�u�WZ�u�WZ�u�WZ�u�WZU�.�Uk����CJ�`��m�	B��QY
+!Ed(�����V\jˍYq�.5eƬ�՗��VZ�U�uZ�U�uZ�U�uZ�U�u]��;��q�.5e�uZ�U�uZ�U�QZU�QZU�QZU�QZU�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U�uZ�U6�bm��۩��Sn�&�LM���u16�bm��۩��Sn�&�LM���u16��Քڲ�VW��5������RmYM�)�e6��Քڲ�VSj��}^����z��W����_W���}^����z��W����_W��l�����}^����z��U�^���W �W �W �W �W*M��;�ʓk�r�mx�6�hM��������r�*mxez�G^����N����mx6� �I���/��������:ܗ������?�����<�a�l�j� ����|B�P�"j�[ej5�|<ġ�Hr$�]�����O1� !�`���yԅ���:@T�Q����5���mt͡�zF1�ӵ3�r�K!��bN�~��V�ƭ�?�[����j����ɯ�&�s���β�r�J��q+:v�bzF1e�6���1�OI�]2�ֽ%�t�Tк� ��]!�E�����bRI�%$����@�w�
�6�Z<�+G��tkX�m��mc���x�6����Z�?�W��u���6�j��'ɴ�bm&��^7]�6��x�q�	�⃹|��^-���N5�|��_9;��N��\��W9���mr���W>�����㛹x��+�GΠ��Pg����ҫ4��M*�J�ҫ4��M*�J�ҫ4��M*�J�ҫ4��M*�J�ҫ4��M*�J�ҫ4��M*�J�>u=��Oc�S����ҫ4��Mr���W>���f����:���S�\�rk�NMs�ɮu95Χ&����:���S�\�rk�NMs�ɮu95��f�X��+��c�\�vk���r�ٮV;4��֕��Һ�ZWS�J�}i]O�+���u>��O��S����>u>��O��S����>u>��Nc���D�Һ��WR�\�Nk����bp�\�!W-�U�br؅\�!W-�U�br؅\�!W-�U�br؅\�!W-�U�br؅X�!V'U��bp�X�!V'U��bp�|�>_(�����|�>_(�����|�/�c��L|�i���1���>_4���J�l����J�l����J�l����J�l���ȅ|���aE�d(�l��m��M�>I�G�6�J�Li\)�+�1�p�4�ƕҸSW
cJ�?iRg�+�1�p�4�ƕҸSW
c��~�x�4������
$�D�`(�P
$�W[e�p�4���M�>I�B���Qx�
/#�t|�n��m��M�>I�G�6��&�8ZaD��Q&�I�j�d^��Ցz�/VE��QY
+!Ed(�����ҫ-*�ҫ-*�>WG���]+��t|�����>WG���]+��t|������+�r��+�r��+�r��+�r��+�r��+�r��+�r��+�r��<O;�+�.��E���#qB�XQY
+!Ed(�����VB�ˍYq�.5eƬ�՗��V\j�\�Ϋ\�Ϋ\�Ϋ\�Ϋ�\�r��5eƬ�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\�Ϋ\��LM���u16�bm��۩��Sn�&�LM���u16�bm��۩��Sn�/U�^���VSj��\Ʊ|�l�D�$�/U�^���W1z�b�\�깋�s���}^����z��W����_W���}^����z��W����_W��l�����}^����z��U�^���W �W �_"M��/W���Bm|Л_4/W���5K������X�J�//Reש2�bLSX��I�/\!��7��M�p�k/�������:ܛg��l�Pm�*CŦ�<ZmB0��F��ƫPn�+J�A1���Z��י�H Z�ĢHr$����~X^M��p7��I�yԅ�����4鎦�]:��t�kޑ�jzF1�ӵ3�r�K*��4����ߣ�M�G�Ib�q%�qĖߡ�-�C�[~�$��I��8����KC�5�G�j�1Ư��)�-������9jf �Ö�jGSj�M{�Q��Lo�םd.��&�CX������bRI�%<�e��@�z��&���V�5�kl�##ڇ�Cl�*m�%Mc���x�/_��[U�u�W���M16�Lw$�n�M6�PM�k�r�mܼ[w/�kŴ��m6�[w/����'��ƾvq���k�gr��ܼsk�ϡE�QD��_knMr���W>���ֹ\��+�Z�s�\�}k�ϭ*�J�ҫ4��M*�J�ҫ4��M*�J�ҫ4��M*�J�ҫ4��C�S�J�ҫ4��Mr���W>������Ƭ[q��jŷ�mƬ[q��jŷ�mƬ[q��jŷ�mƬ[q��jŷ�mƮsq���j�7��Ʈsq���j�7�ͮV;5��f�X��+��c�\�vk���r�٥V;4��f�X�ҫ�Uc�J�viU��*�٥u94��&����+��bs\�Nq���Urx�\�!W-�U�br؅\�!W-�U�br�Q|�_'��E�pQ|�_'��E�pQ\�W'���ErxQ\�W'���Erx�|�>_(�����|�>_(����J�l����J�l����J�l����J�l����J�l����J�l����J�l����J�l����Qx�
/#�t|�n��m֕ҸSW
c\�?k�g�s���u��γ���~�:���Y�\�>k�'�s���u��γ���~�:���Y���~�x�4������
$��L|�l4���\�?k�g�+�1�p�4���M�>I�G�6�J�Li\)�+�1�p�4�ƕҸSW
`���8[�`|�lՑz�/VE�ȽY�!Ed(�����>WG��\����\�����]+��t|�����>WG���]+��t|�����>WG��\����\����\����\����\����\����\����\����J�bm֩��\,HE�+X�<�<��P��VB��QY
+!Ed(�����V\jˍYq�.5eƬ�՗��V\jˍYq�.5eƬ�՗r���sjˍYk�V��k�V��k�V��k�V��k�V��k�V��q��V1Ƭc�X���5cj�8Ռq��V1Ƭc�X���5cj�8Ռq�.5eƬ�՗��V\jˍYq�.5eƬ�՗��V\jˍYM���u16�bm��۩��Sn�&�LM���u16�bm��۩��Sn�&�Lk�/W����WSj��}k��&����_W���}^����z��Wֱyk��yk��yk��yk��yk��yk��yk��yk��yk��yk��|�X�A6�A6�A6�D�_"^�������z�<�_%^�5�4�bM+X�J�8N/\&W�-c�cX��8_�ge�M�p�k/���ٶu�6ηf����?��g�{P�Pj-1���<g�cl�?m�'�c�ݶF6��B�L@�#>�A�Ё�%:C�&�C_���p7����u#�QԂ�pM:c��N���6���ƧN����q4�-�������1�cH~&�qĖ���8i�n��B�锅��)w�R�L�߯LD߯LD߯LD����JJ�&?�����P�����������n&�帖_ьwLck�mk�:��L���޷���o�;|�<�G�"�y�.�)��-�1)��+G����l�$m��֠u�F���P�<J�g�SX�-k&���m��^�O׮�ۅ��p�W�6��&�M�k���A6�PM�k�r�=ܾOw/�k�'��ƾrk���r�ٮ_;4�����X	�_;;�nN5�|��_;8���5�|��_;8���r���W>���ֹ\��+�Z�s�\�}k�ϭr�ٮV;5��f�X��+��c�\�vk���+���u>���f�X��+�j�7��Ʈsq���j���9ƮNq���j���9ƮNq���j���9ƮNq���j���9ƮNq���k�'��ƾrq���k�'��ƾrk��mr�ͮW9���6�\��+���s�\�sk��mr�ͮW9���6�\��+���b�\�[i]NMr�m�V-��ŷ�=ƮOq�����J�O
+���<(�O
+���<|�P/�����@|�P/�����@|�P/�����@|�P/�����A�^6U�a�^6U�a�^6U�a�^6U�a�I�Z�u�I�Z�u�I�Z�u�I�Z�u�^6ZU�e�^6ZU�e�^6ZU�e�^6ZU�d|�n��m��M�ҸSW
cJ�Lk�g�s���u��γ���~�:���Y�\�?k�g�s���p�5���|�8O��Y�\�?k�g�s����>k�g�+��>p����J�l����\�n����s���u��γ��ҸSW
`�&�k�g�s���u��γ���~�:���Y�\�?
:�!G[d(�l�m�
�!WD*�]��t|�����>WG���]k�ֹ]k�ֹ]iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�iW�q���_1ƾc�|���5�k�8��q���_1ƾc�|���5�k�8��	��bB�/��r�nc-�hp��a����]+��t|������+��s��;��w+��W1ܮc�\�r��5eƬ�՗��V\jˍYq�.�s��8՗��:�s��:�s��V\jˍYq�.5eƬ�՗��V1Ƭc�X���5cj�8Ռq��V1Ƭc�X���5cj�8Ռq��V\jˍYq�.5eƬ�՗��V\jˍYq�.5eƬ�՗��V �V �V �V �V �V �V �V �V �V �V �V �V �V �V �W1�I��^W��m]M�����^Z��z��W����_W���}^�����^Z��^Z��^Z��^Z��^Z��^Z��^Z��^Z��^Z��^Z��_ �/�M��M��^�/W���憱xyz�<�$ҵ�Íb��l�2�8N6��C��X�.�:��gZ;l�~j`�X����:�[g[�P�sj�mC�ɶ���� x6�̌n��� 9�l�?k�0��F6��B�L@�#y��1(y��7��K ��]y��$.��wNu7Θ�o^�h::f�ֺv�ڇ-Ĳ���ru������5C�5�C�[��n��O�-��_���_����+���-��4[��h�W��n������M���J�8!!Ąߣ�I^�ķ�?�[�&��j�N���:�����_ьwLck�mk�mh�����4���'I�R7���!�������h��$ Z5������ 㭰8�P�(jC���x�5���ݶ������M16�l���X�l�Rm��M��I�k��M��^(&׊	�⃹x��^-���n��ۍ|��/��Us�x�p��]i�5��X	ܼsw/���7r��ܼsw/���7r��ƾvq���k�g��ƾvq���k�g��Ʈsq���j�7��Ʈsq���j�7�ͮV;5��f�X��W9���n��|��_98���5rs�\��W'8���5rs�\��W'8���5rs�\��W'8���5rs�\��W'8��N5�|��_98��N5�|��_98��N5�|��_98��N5�|��_98��N5�|��_98��N5�\��W'5�Ŷ�X��W'8�����|��_(5����@|�P/�����@|�P/����x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���x�iW���&�k�mֹ&�k�mֹ&�k�mֹ&�k�mֹ&�k�mֹ&�k�mֹ&�k�mֹ&�k�m֕ҸSW
cJ�Lk�g�s����>q�Ϛ�Y�\�?k�g�s���u��γ���~�:���	�\�>k�'�s���u��γ���~�:��o���~Һ�-+��Һ�-+���?ۮ7�c��|��8���7��\�?k�g�+�1�p�5γ���~�:���Y�\�?k�g�s���u��������>�G���]��tB��U�
�>WG��J�cJ�cJ�cJ�c�|���5�k�4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��8��q���_1ƾc�|���5�k�8��q���_1ƾc�|���5�k�6���r���нp�k��H���;��;��;��;��;��;��;��;��;��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��V\j�\�Ϋ\�Ϋ�Yq�.5eƬ�՗��V\j˹\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮb�\�깋�s��/U�^���W1z�b�\�깋�s��/U�^���W1z�cl�cl��W����WW���}k��yk��yk��yk��yk��yk��yk��yk��yk��yk��yk��yk��yk��yk��|�X�A6�A6�A6�D�_"^�������*�|��^k����&e�u�ke��Yv�֎�:��gZ;P��:�6�������:ݚ���X�rm��m��m���Ŧ�<Zb�e�x�H��1� F5Z�r֠�@P�+H��7�h:�-��(�����!˽����E�.�\ꎧ@�L��9�׺s�Lck�jgp帖C��iGYY^��1n8���q' ��߯L����[��k��%}|��x
��8��>;+�|vW��쯡��_C㲾��an��~hJ��-��4iAq�-��鈅��)+���ߣ��^��5zc�_��b[�eӵ3��1�E�p:7��, ���Y:O:����"������h Z�C�m�V�[ej5�#��6��P�<
g�SX�0k&׋Uz�?^�O׮��m��M�[.�Mz�i�Rm5�M��I�ש6�mx��^(&׊��{�x��:�k�&�\��:���`�>^�Ӆ� �5㛍x��^9�׎n5㛍x��^9�׎n5㛍x��^9�׎n5㛍x��^9�׎n5�|��_98��N5�|��_98��Mr�ͮW9���6�\��_98��N��۹x��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��W'8���5rs�\��W'8���5rs�\�ү�U�J�riW�M*�9�_'4���|�ү��U�sJ�Ok��r�A�_(8׍��ү*�ү*�ү*�ү*�ү*�ү*�ү*�ү*�ү-*�ү-*�ү-*�ү-*��$ۭrM��$ۭrM��$ۭrM��$ۭrM�ҸSW
cJ�Li\)�+�1�p�4�ƕ>I�G�6��&�$ۣ�t|�n��m��M�Ҥ��T��\�>k�'�s����j��mW���u�\n�����q�ڮ7[U��j��mW���u�\n�����q�ڮ7[U��j����7��\�?k�g�+�1�p�4���\�n��)������w<Z�7���|��5γ���~�:��o������>q�Ϝo������>q�χ������?ۣ��tB��U�
�!WD*�]+��u�_1�_1�_1�_1ƾc�|���5�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�k�8��q���_1ƾc�|���5�k�8��q���_1ƾc�|���5�����#���pQE:���&�Yw/w/w/w/w/w/w/w/w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1Ƭ�Ֆ��k�V��k�W��V\jˍYq�.5eƬ�՗r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�깋�s��/U�^���W1z�b�\�깋�s��/U�^���W1z�b�}j,m�v�y^���u6��Wֱyk��yk��yk��yk��ym�v�'m�v�'m�v�'m�v�'m�v�'m�v�'m�v�'m�v�'m�lm�lm���e�%���x�z�\�^.k�������+X�8�/5�Í�L�l�.�:˵����u���MC�3P� �:�6η֡���?�ڇ��l�[m��m��m�x�-1Ŧ x6D���?t���09�̌-y�2�L@�#y����rHXG���!��C�{!�� ��]y��$.�V.�GR��4�6����N����q,�-�������1�o�&� ���C�c~�1����_�U������5��hnKhnKhnU�hnK\Y���ܖ(��W���W���|��د����_9\[��}|����O����~)+������j�1�o��+'Y�9n%�N���pkK�tTv�������:O:����.���-�2���- �B��6�>�ej5�V�Z�qטt@�j�ĩ�x�5��ֱ�`�p�/\'��	����M�[)�ez�i�Rm6���^��kԛaz�l&׊	��mx��_'����m&��_9<������(�P�lG�rM�ܓrw$ܝ�7'rM�ܓrw$ܝ�7'��Ƽsq��k�7��Ƽsq��k�7��ƾrq���k�'��ƾrq���k�&�\��+���s��|��_9;��n��۹x��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��_'������{�|��$����\�[k�kmr�=�^'�����x�ү��U�s\�Pk��r�AƼl8׍��ү*�ү*�ү*�ү*�ү*�ү*�ү*�ү*�ү-*�ү-*�ү-*�ү-*��$ۭrM��$ۭrM��$ۭrM��$ۭrM�ҸSW
cJ�Li\)�+�1�p�4�ƕ>I�G�6��&�$ۣ�t|�n��m��M��8O��	�\�>k�'�7[U��j��mWs����j��mW���u�\n�����q�ڮ7[U��j��mW���u�\n�����q�Ϝo���~�:��W
cJ�Li]m����w<���sŪ�x�]����|��8���s���u�����7���|��8���7���|��4�ƕ�ҼSW�`�}���B��W�
�>_G���}/���|����\����\������>_G���}/���|��ֹ'M��5�M�1�z�\�p��^\k�}q��5�ƾ�����_]�˹yw/.��ܼ���r��^]�˹yw/.��ܼ���r��^Si6&�l^�Pkh��Z%��M�����}w/���ܾ���r��_\j�]q��5uƮ�����W\j�]q��5uƮ�����W\j�]q��5uƮ�����W\jˍYq�.5eƬ�՗��V\jˍYq�.5eƬ�՗��V]��}w/���ܾ���r��_]��}w/���ܾ���r��_Z��^Z��^Z��^Z��^Z��^Z��^Z��^Z��^Z��I�ĝ�I�ĝ�I�ĝ�I�g�p�g�p�g�p�g�p�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�gZ&�©�p�6����y�u�:̈fZ�	v��\@� u�:��g����)��j⚇����@� �<@5MC�P�vy�o3�m�x�	��`@�l<�ƛ��l���1�x�H����7t�ʝ r��Z&����rH��D�؁h@�D� �԰�� �����uGS�&�t�S|��A�Ӷ��Ӷ���Ơ帖_��Vo������0[�2��D'��CH?	p����������^�1b�ʾ5xjM��5&�^�n��I�W��J��I�W��J��I�W��J��B�_E�[���|�������-��_�E���!h�߯L�4��b��o�~������sK�1�OH�5:f�ڋ�S^X7����ł��7�*��!��b����bSըZ6ρ��ZH�+I
�h�Z�j�[daP�"k�c��z�7k&c�ݶ�[g�U��Z�Y�X�Lk��[uz�n��-�ۅ��p�]�6����w8[�a��l;�-�MA��Nk�kmrMm�I����n��۹x��^-���n��۹x��^-��iɴ�rm&��I�&�iɴ�rm&��I�5��6�\��_9;��i��sX�Pm�����w/��ŷr�mܼ[w/��ŷr�mܼ[q��k�Íx�q�5�aƼl8׍���I���6��&�w$�n�Mܓi��m7rM��u���ù��w8[4���&��I�5���MAƓPq��i5MAƓPq��i5�x��/���{\�Ok���r�=�_(5���9�_(/]m���~�<M��Y�x�k��6�x�iW���x�iW���x�iW���x�iW���&�k�m6�&�k�m6�&�k�m6�&�k�m7�1��Lq�Sn��1��Lq�Sn��1��Lq�Sn��1��Lq�Snƹ�|�8O��	�\�>k�'�s���p�5���|�8O��	�\�>k�'�s���p�5���|�8O��	�\�>q�ڮ7[U��j����7[U��j��mW���u�\n�����q�ڭ+�ݥu�����J�j����J�j����J�j�����|ҿϚW��J�>i_��+����5�v��n�<M�牻\�7k�&�s�ݮx�����J�j����J�j����J�j����J�>i^)�+�1�x�4����^B��Qy
/!E�^ZU�^ZU�^ZU�ƾ�����_ZU�^ZU�^ZU�^ZU�^B��J���h/^+�ǂ�����ƕyq��5�ƾ�����_\k�}w/.��ܼ���r��^]�˹yw/.��ܼ���r��^]�˹yw/)������i6;��r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r���s��;��w+��W1ܮc�\�r���s��;��w+��W1ܮc�\�r��_]��}w/���ܾ���r��_]��}w/���ܾ��ֱyk��yk��yk��yk��&��&��&��&��&��&��&��'k��'kv�'kv�'kv�'m�6��m�6��m�6��m�6�'j,j,j(55��
C��C���ơP�cP�A�p��p��8Pm�*�g
�����:�5���Q�ȁ�e�p�:�c��3�S���?�/�C�SP� �?�5MC�P�vj��3�m�x-�	��x���y��7���y����~�<�g����j����9S�T�+D�`r&��o��J -BHr$��k����o�;����2��zM�d��A�Ӷ����פc��S;�-�үLr���b�锟4Z!u~|��W���_b���b�e��T���T�N�,��H�0jX�E�c��Z�0jX�E�c�N�$F�FH�+iq+�Rm�4\5�h�܋p�L����4��=�C�������O�q'?�����P�)�#��ڙ��ƧL�R����ޖ
;|���'H��y�o'H��y�OQ��Z5���ZH�+F�
�kP:�#ڇ�l�k��Y�X�-k&C����[g�U�u�5��Ʊ���u�W������M�[)�e6�l��m7s���p��ù��w8[7
s��$���۹x��^-���n��۹x��^-���n���m&��I�&�iɴ�rm&��I�&�iɴ�s\�sq���k�'r�mz�Okjc�A���ŷr�mܼ[w/��ŷr�mܼ[w/��k�Íx�q�5�aƼl8׍���^6�6��&�w$�n�Mܓi��m7rM��I��n��m��w8[�aƓPq��i5MAƓPq��i5MAƓPq��i5MAƓPq��i5MAƓPq��k�Íx�iU��5�az�n������kg���uƾl����J�l4���J�l4���J�l4���J�l5�6�\�i��6�\�i��6�\�i��6�\�i��)�7
c��p�8�)�7
c��p�;�g��Y���~�u���g��Y���~�u�����|�8O��	�\�>k�'�s���p�5���|�8O��	�\�>k�'�s���p�5���|�8O�n�����q�ڮ�����n�u�\n�����q�ڮ7[U��j��mW��Һ��WY�J�j����J�j����J�j����J�>i_��+����4����|ҿϚW��\�7k�&�s�ݮx���v��n�<M�牻J�j����J�j����J�j����J�j����J�>i^)�+�1�x����^B��Qy
/-*�ү-*�ү-*�ү.5�ƾ����ү-*�ү-*�ү-*�ү-*�WG������m����A�I�U�ܼ���r��^]�˹yw/.��ܼ���r��^]�˹yw/.��6��ה��^Sk�myM�)��ܾ�ו�M�ԛ�6/RlM�.��6��ה��^Sk�myM�)��ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��^Z��^Z��^Z��^Z��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d��I�d�@�D u�8Uh�BZ!�P�ֈ@�T u�8Uh�BZ!�P�©�u�5��C��P�< u�:̵�X��`��1�u���MC�0�� @�  �?��m���x�j������� x�	��x���<3���</3���x���I�t��V��-t�ʛ����V��J�7IZF�-�P�`Jy��o2���]�E�.�\�Χo�U���N��o];hkC���ڙ�9jf 帚_��SW��,i$'�zau|W�%}|��}Ϛ.��hY��iR�2��,`"�[_&��f����ߛЬo��V7��+�z���
��ޅc~oB��7P����i�Z��"��J��I�W�������C�@�|���W�����O�q)#�1���帚];S1=&�wt�1�]:���p:7���t�v�@Cp.������1)� Z��&��6�+F�eh؀��F#Zǁ��&�?���kX�-k&c��z�7m��V���kg�c���u�5�����z�?^�O�n�m��M�[)�e6�l��m7s���p�i5MAƓPM�ӓi4��M96�NM�ӓi4��M96�NM�ӓi4��M96�NM�ӓi4��M96�Nq���j��r�=6�P^��c���8Zm����^(&׊	��mx��^(&׊	��mx��I���6��&�w$�n�Mܓi��m7rM��p�Sn�m��M�[)�e6�l��-�ۅ��u��n�����w8[�aƓPq��i5s���p��ù��w8[�a��l;�-��&�Ҥ�T��J�PiW���x�iW���x�/�U�a��?^�Z�׋U6�>q�S�u�I�Z�u�I�Z�u�I�Z�u�I�Z�u��Lq�Sn��1��Lq�Sn��1��Lq�Sn��1��Lq�Sn��1��?w:��γ�s����?w:��γ�s���p�5���|�8O��	�\�>k�'�s���p�5���|�8O��	�\�>k�'�s���p�Z�U�p�\n�w����0w?���s����0w?���s����0w?�����`�?����\�0k��s���x���v��n�<M��U�x�Z�U�x�Z�U�x�Z牻\�7k�&�s�ݮx���v��n�<M�牻\�7k�&�s�ݮx���v��n�<M�W�U�x5ZW�U�x5B��Qy
/!E�(����yiW��yiW��yiW���_\k�}iW��yiW��yiW��yiW��y
+����I�n8�,q�X�$�*��^]�˹yw/.��ܼ���r�I�6�bm&��M���i6&�lM�ؽI�z�b�&��M�ԛ�6/Rl^���W]��my^�ؽI�6������^Sk�myM�)��6��ה���_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��_]��}w/���ܾ���r��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה���$�N�$�N�$�N�$�N�$�N�$�N�$�N�$�N�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8Py�m3���u�<ζ�����:�g[C��hy�m3���u�<ζ�����:�g[C��hjg��Y��(�����y�����XǙ���?�ڇ����@�  �y�/o3���x�y� ���!��@�s<\�g����[<�db�̌i��ƛ��n�H����?t����ݿ����ai`T�ե����V�������$o�tr.�@�"S��%=K�]��*��(�Au�&�1�޺v�ֽ#���r�K/��++���G�X�	���������>4+�|vW��f��B�^��i�d���M��� �Bj'�=
"ă��/^$�,H1x-�c�[ ��A���i1l����
�m	�:�+�u"X�2�_���ʾ���H?	?��"W��	�$�������f'N�K/H�5�Q��nF��N�Τy�)'H��y�o'H��y�OQ��|	�2�m�V���kl�kM��M�x������T�<Lǉ�l�7m��V���m��V���kg�c���u�/\'��	����^�۫�[uz�n��m4ۭ��u���ù��w8[	��m&��I�&�iɴ�rm&��I�&�i��
z��p��\)��
z��p��\)���{�|��^(&׊ԛaz�l5��X�i�׊	��mx��^(&׊	��mx��^(&�-�ۅ��p�Sn�m��M�[)�e6�l��-�ۅ��p�Sn�m��M�[)�e6�l��m4ۭ��u���ù��w8[4���&��u��n��m��M��i�[M6�i��m4ۭ��8[s���8[s���$�mrM��$�mrM�үrM��u����ɷ��m�|�u���)�7
c��p�8�)�7
c��p�8�)�7
c��p�8�)�7
c��p�8�)��Y���~�u���g��Y���~�u���g��Y���~�u���g��Y���~�u���g�7[U��j��mW���u�\n�����q�ڮ7[U��j��mW���u�\n�����q�ڭs���u���f�7Y���`��;�������`��;�������`��;�����\�0k��s����5����`�<M�牻\�7k�&�sŪ�<Z�sŪ�<Z�sŪ�<Z�7����`�x8�7����`�x8�s�ݮx���v��n�<M�牻\�7k�&�+��Ҽ�+��Ҽ��|���q�N>I��;\���;\���;\���;�yw/.��ܼ��;\���;\���;\���;\������ү-rN�$�rN�$�rN�^]�˹yw/.��ܼ���r�I�6�bm&��M���i6&�lM�ؽI�z�b�&��M�ԛ�6/Rl^���W]��my^�ؽI�6������^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה���$�N�$�N�$�N�$�N�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X�8X u� u� u� u� u� u� u� u�t��'ZWI֕�u�t�i]'ZWI֕�u�t�i]'ZWI֕�u�t�i]'ZWI֕�u�:̈f^g�w��\@�.�<F<��w����<_�'���� @� �<^�g�ۤ�}t��C���� x��.o3�m�x-���=�F4�dcM�F7]$cu�x�H��I�t��R���*o�҆��(,B�Ќ�Z#K�5������y��`9y���p= *��7���N��;hk];SmC��jGY��ef�ɣH~%�!Ą��L.����^�Ӌ�b��|��ԜJ��R%�o�:�o��Vd �o�F�o�x��<[��-���������������y�ߘU�-�b�1��qc�E�i�,�8Yj4�Gb�uxjF�}�I���'��h.߯L�ߣ�9^�$��)�#������]m�`����޷�*��y��Χ]1� �ځ���%=^e���$����b5�x��&��D�<J�g�Sl�*k&c���x�6��v��n�?��g��l�7m���c���u�5�������/]m�뭺�u�Sn�m��M�[.�a��l;�-�s���p��ù��w8[�a��l;�-�s���p��ù��w8[�aƓPw8[�a��l;�-�s���u��n�����w8[�a��l;�-�s���p������^�۫�[uz�n�]m�뭺�u�W���m��M�[)�e6�l��-�ۅ��p�Sn����^�۩�e6�l��-�rM��I���6����^�۫�[uz�n�]m�뭺�u�W�����q��n7[M��i��-����p�\n�\�n��)��Y���~��&��ɷ���~�u���g��Y���~�u���g��Y���~�u���g��Y���~�u���g��Y���~�p�;�'��	��|�p�;�'��	��|�u�Sn��m��M�ک�[U6�j��mTۭ��u�ZW�U��ZW�U��ZW�U��ZW�U��ZW�U��ZW�U��ZW�U��ZW�U��7q���n�ws����0w?�o��ĵ��0w?���s����0w?���s����5����`�?����\�0k�&�s�ݮx���v��n�<M��U�x�Z�U�x�\o����0q�o����0q�牻\�7k�&�s�ݮx���v��n�<M�W�U�x5ZW�U�x5G�8�'$��|���v�'k�v�'k�v�'k�wr��^]�˹yk�v�'k�v�'k�v�'k�v�'k�v�'k�v�'k�w��7δi6&�lM�؛I�6�bm&��M���i6&�lM�؛I�6�bm&��M����6/Rl^�ؽI�z�b�&��M�ԛ��my^�ؽI�z�b�&����_W�6/Rl^�ؽI�z�b�&��M�ԛk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^Sk�myM�)��6��ה��^W�6/Rl^�ؽI�z�b�&��M�ԛ�6/Rl^�ؽI�z�b�&��M���I�d��I�d��I�d��I�d��p��p��p��p��p��p��p��p�@�@@�@@�@@�@@�@@�@@�@@�A�x�t�+�'��I��x�t�+�'��I⩿��7�����8�������o����q���7�����8�������o����q��y���g�wI�1�x�t���S���<_���3��{y�/n�����<]'���� x>��'����#�$bp��� x'�@�H��#��1�F7�v�7o���괠]V��1uhD.��1(t]%����$�oWL�3��Hn�t��t�:I�(�GN�פ����5�Ɍm[��^��zc���S|���-ޙI�^�]^�z��a���ԍe�Ԕ���\J�-F��i0ud �,H1xX���ߐ<�pB�����;��v�b�k~1z���Zߌ^�,H����y�X�����U&ߘ�|-�B��B��B��0�H���xX�Gb������a����H?	7����)'�NW��49�n���]1�jN���nB�Go��o�U���� ���!��7x���t�OW�h�+D�`q� 9#P�F���6��D�<�g�Sl�*m�%Mc���x�5��n�<L���P�0m������?ڭc���u�5��Ʊ���?���b���^�۩�e6�l��m4ۭ��u��n��m��M��i�[M6�i��-�s���p��ù��w8[�a��l&�m4ۭ��u��n�����w8[�a��l&�m4ۭ��u��n��m��M��i�[M6�i�]m�뭺�u�W������^�۫�[uz�n�]m�뭺�u�W������^�۫�[uz�n�]m�뭺�u�Sn�m��M�[.�Mܓi�]m�뭺�u�W������^�۫�[uz�n���s����]��˹��w:ۮ�[u��n��g��Y���~�u���g���m�|�x�]γ�s����?w:��γ�s����?w:��o�����6�>M�ϓo�����6�>M�ϝ��s����>w8O���s����>w8O�n��m��M�ک�[U6�j��mTۭ��u�]��v��n�<M�牻\�7k�&�s�ݮx���v��n�<M�牻\�7k�&�s�ݮx���f�7Y���`��;��	��jm�Z�x���%���jm�Z�x���%���jm�Z�x���%�7�k��Z�x���%�7�k��`�x8�7����`�x8��7����n�x��7����`�x8�7����`�x8�7����`�x8�7����`�x5��v�n�#��a���8c�|Ꮬ1��$�rN�$�rN�$�rN�I��;�'w$�rN�$�rN�$�rN�$�rN�$�7���;\���;��M��M��M�i�6��4ۆ�p�nm�^�ؽu�z�b���뭋�[��/]lklklklklklklklklM����u��u��u��u�z��u놽p׮��^�k�z�\4�N�I�i:m'M�鴝6���t�N�I�i:m'M�鴝6���t�N�I�i:m'M�鴝6���t��^Sk�myM�)��6��ה��^Sk�myM�)��6��ו놽p׮��^�k�z�\5놽p׮��^�k�z�\6��ơ�jv��jv��jv��jv��jv��jv��jv��Ǚ����y��g������y��g����ho����ho����ho����ho����d�x�,#����0�x�,#����0�x�,#����0�x�,#�Ǚ�]�x�y�#g��I�)�x�t�/����xy��g�ۤ��<[�1ٿ���1��x9<�'����#�$bs��Ny��21A��[��1����0������sr�Z`X+L��`�V�b�Ѝ�-�H�H�#Θr<.�@ސE���p:`���\H
�zM�d�GGN�פcC��jGY��G�~��Q�?E��)>h�BW�~W���4��[Z���6Ұ|�o�:�|�M�����[ ��~@����;�a��^F�h�#�r�#�r�#\CW��!�����k�j�5�5y���������~1;~Az1� y�X��������U|ߘA���� ���x4�G�5#[����H?	u~"|�h�4��9��W�c�^�S;��3ZX6����Ӥ��ł��t�u;y��E���O1�����)��- ��! 9#P�F����F�<���l�*m�%M����x�5���` x��C���x�5��n�?ڭ����?ڭ����?���cX�L^�۫�[uz�n�_������W������^��+��ez�l��m4ۭ��u��n��m��M��i�[M6�i�_�ۭ��u��n��m��w8[�a��l/_������W������^��+��ez�l���Ʊ�|�:Ϛ�Y�X�>kg�c���u�/\'��	���~�p��\'��	���~�p��]m�뭺�u�W���m��M�[.�Mܓi���Ʊ���?���cX�Lk�c�1��;��s���u�]ζ���w:ۮ�[u��n�����Y���~�p�;�g�����n�<Lo�����6�>M�ϓo�����6�>M�ϗ�����^�Z�׋Uz�j�^-U�Ū�x�Sn��m��M�ک�[U6�j��mTۭ��u�Sn��m��M�ک�[U6�j��mTۭ��u�]��v��n�<M�牻\�7k�&�s�ݮx���v��n�<M�牻\�7k�&�s�ݮx���f������`��&�%���jm�Z�x&�%���jm�Z�x���%���jm�Z�x���%�sĵ�x���ֹ�Z�<KZ�k\�-k�s���x5���`�<�a�\�7q�\h��0�ƌ-q�\h��0�ƌ-k�s���x5���`�<灃\�0k���r0ݮF���v��i]v��i]v��i]w��p�n��q�n7���4ۆ�p�n��q�n7���7��p�ζ;�lq�mrN�p�ζ&��/^(�nm�M�i�6��4ۆ�p׮�/]l^�ؽu�z�b���뭋�[�[�[�[�[�[�[�[�[���klm��6���]z�\5놽p׮��^�k�z�\5놽p׮��^�k�z�\5놽p׮��^�k�z�\5놽p׮��^�k�z�\5�M�ԛ�6/Rl^�ؽI�z�b�&��M�ԛ�6/\5�M��z�b��^�k��I׮l��\6�'^�m�N�p�d�z��:��m�v��jv��jv��jv��jv��j,jv��ơ�ơ�ơ�ơ�ơ�Ǚ����y��g������y��g��t+FQ�[�0Ⱥ�2�ц[�0�Fo�v��G^"���]x�o�qu�)���׈���G^"���]x�o�qu�)���'�;���?��'��I�)�x�7��g���x����I�	�x>��c�F;7�����ry�O3�m�F':H��I��ъ21A�F4��:cLo���������i�`�0,���L]Z�B7LJzD�GL9tÑ��r<.�@�ם���p:`��]��b����Ә�{�1�������q5+�үG�����q&�h�B���������رF�䱚���
3�[@�Ql�������8K/�4V�fk�O컈m�a�ם��
߁zo��n�m��m�7�M���*�����g�����4���4�QZߐ^�,H�����ߘ�|���[Bi�|�*��T��.)���+��~h|��$-����^�I^�$�Nc���S;����N�������E����U�`�� ��������-�)��- ��'�x@H�#���u�x��&��&�<J�g�SX�0k&c��@�-<D֡�`�<L���l�j����l�j����l�?k�c�1��/]m�뭺��W������^��+��ez�l�_�����u��n��m��M��i�[M6�i��m4ۭ���W������M��i�e��l;�m7s���u�W������^��+�[uz�l�]m�뭺�:Ϛ�Y�X�>kg�c���u�5����|�p��\'��	���~�p��\'��	���~�?�������^�۩�e6�l��-�rM��?���cX�Lk�c�1��5��Ʊ����&�鉷�bm����&�鉷��m�|��;�g��Y���u��������X�0M�ϓo�����6�>M�ϓo�����6�>^�Z�׋Uz�j�^-U�Ū�x�W�����M�ک�[U6�j��mTۭ��u�Sn��m��M�ک�[U6�j��mTۭ��u�Sn��m��w?��牻\�7k�&�s�ݮx���v��n�<M�牻\�7k�&�s�ݮx���v��n��;�������`�x���%�ׁR��T�x���%���jm�Z�x���%���k��Z�x���ֹ�Z�<KZ�k\�-k�%�sĵ�x5���`�<灃\�0k���r0�ƌ-q�\h��0�ƌ-q�\h��0��x5���`�<灃\�0k�s���F���v�n�#���������������������������������w:��p�n��k�v�'k�v�yq�n7���7��p�n��^����z��_����ׯ���^����z��_����ׯ���^�ؽu�z�b���뭋�[����^����z��_����ׯ���M�i�6��4ۆ�p׮��M�鴝�^Z��^Z��^Z��6���t�N�I�i:m'M�鴝6���t�N�I�i:m'M�鴝�I��I��I��I��I�d��I�d��p��p��p��uڇ�]�p��u�g�u�l�6��8m���?� x�'���`��t��?� �@�@@�@@�A��y��'��I��x�t�+�'��I��x�t�*�'��I�@�T x�y�3���x4:H�Γ���8X�o�� q��a`1���o��M�)�������x�o��������f��~,!�����x�o��������f��~t�/Γ�Sxy��g�gI�	�xt� ��1��F;<��gI��#�$b�Oo����=���1A�� vä�o���Lt��$a�7o��傴�]|�g���|	��B6��#,	C��(t]%1�t�$.�ċP�!��5���3Βt�:�9n'Nu7��pM:c�[��91����4�#�Y�C�X��J��p+����,Vҥ,`#��0�H��MD��Ь,a��WYbE����v�aG���))�2m�o��7��߀@���y���"����߁�1��<�;�WHizizizq6�4���k�/����U���
�Ɯ �p�@����ӁJ�ԍb�>;+��lA�U�5�^�Hi��?_��Vt�L�����ӷ��Q�N�
�:`��]�������/!t��,/&�J_�KG{��z�O08����F#Z�q��F�#��6��P�<
��@��T x���h��Z x���kl�j����l�j����l�j����l�j������k-ֱ��k-ֱ��k-ֱ��k-ֱ��k-ֱ��k-ֱ��k-ֱ��k-ֱ���?��Y�X�Lkg�c�1�u�5��Ʊ�|�?��Y�X�Lkg�c�1�u�5����|�:Ϛ�Y�X�>kg�c���u�5����|�:Ϛ�Y�X�>kg�c���u�5������6�>M�ϓo�����6�>M�ϓo�����6�>M�ϓo�����6�>M�ϓo�����6�>M�ϓo��ۭ���&�mTۭ����_�������n���_�������n���_�������n���_�������n�<Lǉ�X�0k&c���x�5���`���_�������n���_�������n���_�������n���_�������n�����������n�����������n�����������n�����������n�x8�7����`�x8�7����`�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�x8�7����`�x8�7����`�F�����ak�Z�F�����ak�Z�x8�7����`�?��?�s��s��?��?��?��?��?�s��?�s��?�s��?�s��u���c��q�n7�I�䝮I�n��q�n7���7��pׯ���^����z��_����ׯ���^����z��_����׮�/]l^�ؽu�z�b������ׯ���^����z��_�����nm�M�i�6��5놽p׮��m�v�'m�v�'m�v�'^�k�z�\5놽p׮��^�k�z�\5놽p׮��m�lm�lm�lm�lm�v�'m�v�'j,j,jv��jv��jv��y�w��y�w��y�w��y�w��t��I�t��I�t��I�t��I����������t�+�'��I��x�t�*�'��I���t��'��I�x@�T�<g�C��ht���$a�I�q����q��cF
o��M�)��<����X# ��0`� X# ��0`� �����3xo� �����7��f�������3���<:O N��F;7�c�̌vy��Β1m�F-�H�������������ъ���,��H��խ������$a�>o��傴�]|����L�,m�hF�քe�(t]�K�`CHbB�I���� �԰��0��p�)9��=&К[�i��{�:�O�,�s���᪽	��_��4>4+��lW��f��JX�E�~aԃ��B�����7��-�
1�#J�i�Jq�Cq6��M�#��!`?�e,�̂��߀�^��Qu�eU��Qu���7yf� �������5�S~4ڎX��-�����x8����#I�+ТК@�_$��(�7����T�H\+��~OLD߯L�ߣ�9�egNc]9�ڇ-����s����I�Y�5�`Cp7�ˠ]!��Ȱ��%���|=D
�7�y�j�֡�j�[da�F F����P x�%B�h��Z x���h��Z�?ڭ����?ڭ����?ڭ����?ڭ����?�ǋu�x�Zǋu�x�Zǋu�x�Zǋu�x�Zǋu�x�Zǋu�x�Zǋu�x�Z��cX�>kg�c���u�5����|�:Ϛ�Y�l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j�������^�Z�׋Uz�j�^-U�Ū�x�W�����^�Z�׋Uz�j�^-U�Ū�x�W����n���_�������n���_�������n���_�������n���_�������n���_�������n���_�����X�0k&c���x�5���`�<Lǉ�X�0k&c���x�5���`�<Lǉ�X�0k&c���x�5���`�<Lǉ�m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	�����`�x8�7����`�x8�7���Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak��`�x8�7����`�x8�7���Z�F�����ak�Z�F�����ak��`�x8�7����w<n�����s�������w?��������s��u���c��w?�������w��u�����w��u�n���q��7]z��_����ׯ���^����z��_����ׯ���^����z�b������뭋�[��/_����ׯ���^����z���4ۆ�p�nm�M�k�z�\5놽p׮l���;l���:��^�k�z�\5놽p׮��^�k�z�\5놽p׮l���;l���;l���;l���;P��P��P��P��P��P��P��P��P��P��P��P����D�?�<��O3���T�<U:OM����������)[��+x�o���╿�R�������<$a�I�q���H��0�`�X� �ŀ;����t�����`�X< E��`�X< E��`�X< E��`�X<<� �3�3���<:O M���ю����#�$bۤ�Nt���0:{���+T%j�`�,��H���[����խ���X+O��;U���Ki�`�0_��hTX>�ա`J,	C���.�Q��l]��1'L^w{���0��w��N��o�ь޺s�zM���chrc����bC�M^�$��ze'����.��\S+�RmƜ�|�Y�o��V$�x*�o�!o�Ғ��M������e�n%���~N-b����!��|����*�h,E�Z�~z47�MI�
�2='�����:`����~e�1��j��I���mGx|�ȅ����[A���������m���7*��Mb�\6+��$�E��~�2�~�$�zc�Ö�bt�Sj�Φ�9:�������β,*F�I7 �9p��`9y7�R��Z;�g���V�<��� rA 9#P:����ba�& F	�����P�<
g�Č*y��O20��F5��`�<Mڇ��P�7j&�C�ݨx������~�<O�g��l�?m�'����x������~�<O�g��l�?m�'����x�����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j����l�j�^-U�Ū�x�W�����^�Z�׋Uz�j�^-U�Ū�x�W�����^�Z�׋Uz�j�_�������n���_�������n������`�<Lǉ�X�0k&c���x�&�&	���m�`�x�&�&	���m�`�x�/^�ׁj��Z�x�^�ׁj��Z�x��&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�&�&	���m�`�x�;����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F�����ak�Z�F��7s��x����w<n�������s�������w?��[ζ&�,M�X�x������s��u�n���w?��������s�������^����z��_����ׯ���^����z��_����׮�/\(/\(/\(/\(/]l^�ؽu�z�b��^����z��_����ׯ����뭋�[��/]l^���:��:ؽp׮��^�m�N�$�N�$��z�\5놽p׮��^�k�z�\5놽p׮��^�mC��C��C��C��C��C��C��C��C��:�C��:�C��:�C��:����?� �@�`�����C��:�C��:�C��:�C��:�3���D�<W:O������������0�`�<X<����`�8X<���㤌<�#7�t��e����q��a`�X� �ŀ;����t���c躌}Q���1�]F>����u�.�K�"���x, ��"���x, �$`I�xo�����},݋ w2���F-��t�������%j���Pt���Z�,����o���V�K�a`�L,�傴����Ki�`�0_��hT�E�Љ���P�9F���k�!��L�:`���]0~��S�-�H�Φ����jgG��Z�N��帚���bC��^�$Ѥ����_��4>4+���W���,U`4�f�7�XX�b�i������\9q6��O����+1�2����N�"ߢ�#I��`��B�_4,X���W��b
�|��2�_4,���Z�~��W���@�?e�=5y����P���ka���V�m)(�"�`�C�l�W���B�Z��W�f��B��_9=�+�h�W��n��M�?�_�q4�����S�mk�nG����םdX<�v�I���!�������%���|=]%h���y��b rA� V�^`qטu�"#�$`���t��n�0M�(t�� r�H�@�-<D��@�0<���x������~�<O�g��l�?m�'����x������~�<O�g��l�?m�'�����[g�U��[g�U��[g�U��[g�U�x��v��n�<Mڇ��P�7j&�C�ݨx��v��n�<Mڇ��P�7j&�C�ݨx��v��n�<Mڇ��P�7j&�C�ݬx��v��n�<�ǁ�X�7k�c�ݬx��v��n�<�ǁ�X�7k�c�ݬx�5���`�<Lǉ�X�0k&c���x�����Z�<[g�kl�-m�����z�-^�W�����z�-^�W�����z�-^�W�����z�-^�W�����6�0M�Lo���6�0M�Lo���6�0M�Lo���6�0M�Lo���6�0M�Lo���6�0M�Lo���6�0M�Lo���6�0M�Lo���܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�܌-w#]���r0�6T�*M��&�ʓ`�I�r��9Rl�܌-w#]���r0�6��є�2�FSh�mM�)��6�bm���ŉ��o�o�o�o����o&�,w?��������s�������w?��������&��&��&��&��&��&��&��&��&��&��&��&��&��&��&��5��Mc�X�D�:�5��Mc�X�A���?�k�5����cōcōcōcŋ��z��_����ׯ���^��c��:�c��:�c��:�C��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:�c��:������������������������3���D�?�<��O3���D�?�<��BZZZZZZZZ���S��hy�3�+��8�<:O�����8�<�O.��ˤ�2�<�O��e����a���2X�,� �ŀ;�.�C7�h�� �����;�{o��e�;�`�X� �ŀ;�`�X� �����я����я����я����я����я���X� �e�;�No����9���
��Z�������խ6��i��ku��[���0�|&
��u�|X>���`�7_���-
�ա��"tĢ7LJ#G(�LC$tÑ��C t�8�yǅם�.����p=%$��u�r���hM+֦to��׿��׿��ڿ���4���	�I铅��L|��.���\iڑ��[J̱�$�����5�~@���8�AEk�N�����ho��o���i�L-2���l[�F,E�Bň��@��>g�c����/����>`^�<����(T�|b���lE��4ʽm/�C����L��3<���aqi�m��o;��*ѿ ��ߐX����ЛHX��D�@����&�[��f�|����O�-���KW�YY^�2��1����6�'S^�ۃz逭�� ���<�wL��1$.�\���t����h�- �eh�̭y��b rA� V�^`qטt@�#��10L@�#� � r��T�#
��r֠��-j�Z�r֠��x5��|�<����P�>j�C���x5��|�<����P�>j�C���x��v��n�<�ǁ�X�7k�c�ݶF6���`�#da�l�0m���0��F6���`�#da�l�0m���0��F6���`�#da�l�0m���0��F6���`�#da�l�0m���0��F6���`�#da�l�0m���0��x�����Z�<[g�kl�-m������F5¦�T�#
��aSP�*j�MB0��F5�¦�T�#
��aSX�*k�Mb0�z�-^�W�����z�-^�W�����z�*^�
������z�*^�
������z�*^�
������z�*^�
��������*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*w<
���s����*q�
�o�����*q�
�o���܌(w#
�r0�܌(w#
�r0���*q�
�o���6��є�2�FSh�mM�)��6�bm���ŉ��o�o�o�o��b&��z�Az�Az�A6�bm���ŉ��o&�,M�X�x�6�bm���ŉ��	��	��	��	��	��	��	��	��	��	��	��	��	��	��	��c�X�D�:�5��Mc�X�D�:�5����c����X�A�x��x��x��x��x��x��x��x��x��x��x��x��u��]�u��]�u��]�u��]�u��]�u��]�u��]�u��]�u��]�u��]�u��]�u��]���������������������������������?�<��O3�s��D�?�<��O3�s��D�<U:OΓ�S��\�<U:OΓ�P���x4<������#:O��e����a���2�ц[�0�Fo����]����av��.X�,˖ ���j8��G,ߋ w�L� 镯e���|=�
�E��`�X+A��1uZ�.�\��k���sU�b��]V�� �ŀ;�`�X� �ŀ;�`�X� �ŀ;�`�X���!uZ���Ӌjy`�O,�債@]|6���X>%��X>%��0�|&��uh~.��2Ѫ.���Ѫ.�����Z="Q@��"tĢ7�9zC��LC$t�2G�C t��L�='��逫�L_�`+��(�'N��_�Բ[Bi^�3�~��^�m�r�MM�?���pMW�h�-Ţ`�W�%|�
�4��Ɯ�,`�H����/����^F�h��\9o��6��DYcΘ8eӇ�L��q�~��ث��X�ӿ���0|���J���"�^c��B������M6���|�-��w��`^�<���ث�@i�n|���0~��[�<�;�-A��Ӹ"��J�o�x$<�|��XX���^ �%|m&���I�Ż�'�u~A�1�G�k�n&�z��-�c��mN���(�Lo�0�z@U��y��G.�r�o���Jz�D����t�����V��ςA��+Q�����<��O09�D��<��O2�M�V��¦�T��� �@9kPZ��� �cT@�j��Q1� F5Dƨ��#�cT@�j��Q1� F5Dƨ��#��0��F6���`�#da�l�0m��@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �@9kPZ��� �B0��F5¦�T�#
��aSP�*j�MB0��F5¦�T�#
��aSP�*j�Mb0��F5�¦�T�#
��aSX�*k�Mb0��F5�¦�T�#
��aSX�*k�KׁR��T�x/^KׁR��T�x/^KׁR��T�x/^KׁR��T�x/^N�S��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�I�aBmP�F&х	�aBmP�F&х�S��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�N�aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���mz��A��z���Q��2�x �x �x�^�Q/^+���׊���m�6�D�F"M�;�;�8�,q�X�x���c���Ŏ7�o8�,q�X�x�^�Q/^(��K׊%����z�D�x�^�Q/^(��K׊%����z�D�?�6�������?�g�Cl�\�?�6��ͳ�sl�\�<Q6�M��l�D�<Q6�I��o&�,M�X�<X�<X�<X�<X�ׯ�X뵎�X뵎�X뵎�X�_����ׯ���^����z��_����ׯ���^���������������������x��<Pj(���&�≨x�j(���!�P��@�< x�?�*��������x4<��3���x�y�3�+��J�<R��Ï20�̌8�#�H��0����7�q��)��7�`����т��8��a`1���,��;�.��A��@B���]|>����uZ�.�\��k���sU�B��]V���!uZ�.�\��k���rU�B��]V���!uZ�.�\��k���r,�� w1uZ�.�\��:q`�O,�債<]|6��a��Zm�Z�,����V������|&�C�u�|.��գT]Z5E����Z�e�S�ZB�t�P�DoHr:�#����zA��B$��zO;�Ӂ]�
�zJ;��\IGI:f�zGR�9m	��c7�鸛_�q6����4����|�O�-�4?���W,Q��u`XϒD[Bi��k��bǃ���¼�q�2m�|��e�:`�r�űM�[n,E^��0��8�\o�ƚjۿ�X8eӿ��dW����7�c�̯���gL����������񦚇�E�M�g|�P���>hM�
���/����q|��o쵊;�g�����"������zE��$U���_4hSp���������Hi��?���VGY�^�2�rc];hk]3p:�;z逭���^�b�u8�I�7C%/��)~���2��Z�O�I�@�>	g�#��$y������V��J�7IZF�+H�%i��#t��b r� 9@��@P (��BiŠ-y���20��F���יZ�#^daǩ-y���20��F���יZ�#^dakP�*j�MB0��F5¦�T�#
��aSP�*j�MB0��F5¦�T�#
��aSP�*j�MB0��F5¦�T�#
��aSP�*j�MB0��F5¦�T�#
��aSX�*k�Mb0��F5�¦�T�#
��aSX�*k�Mb0��F5�¦�T�#
��aSX�*k�Mb0��F5�¦�T�#
��aSlP��6���9ClP��6���9ClP��6���9ClP��6���9CX�*k�Mb0��F5�¦�T�#
��aR��T�x/^KׁR��T�x/^KׁR��T�x/^KׁR��T�x/^KׁS��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�N�S�P�F;���aC�P�F;���aC��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S�P�F;���aC�P�F;���aBlM6&�M������`�i�q4�8��P�F;���aB���A��z��FW���^�^�^�Q/^(���׊���r��z�z�6�D�F"M�;�;�;�8�,q�X�x���c���Ŏ7�o/^(��K׊%����z�D�x�^�Q/^(��K׊%����z�D�x�^�W6�������?�g�Cl�hm����sl�\�?�6��ͳ�sl�D�<Q6�M��l�D�x�6�bm���ōcōcōcōcŋ��z����X뵎�X뵎�X�_����ׯ���^����z��_����ׯ���^����z����6��6��6��6��6��6��6��5��C�P�D�<Q5MC�P�\ �?����������x@�<�<:O�����8�<:O�����8�#<�Ï20㤌.�#�H���c���7�`����т��0SF
o��M�(�F
,�
�r��]V�U���p�8u��.�E��躭sU�b��]V����1uZ�.�\��k���rU�B��]V���!uZ�.�\��k���rU�B��]V���"��]V���!uZ�X+S�jy`�O_
��.��Z�,����V��uh~.��ա���?_Ιh�V�Quh�t�B�L�-t�B�L�*IE�r&�DoHr:��h�LF� �����g�y�D����t�W{�Q�OIGy:`+��\ꎧzGR�9m	��c7��Sk_�SmU�i��_^�1^�	_U��__9=_b��ӁCNo&�|�Uxߐ^�q�Z+���țnL����.�?�i6�l�:X��,`�b�w+�o��?�W�Ӗ>o�4�2�����w�b�K�ݿ
�+�|������o����/���zO��o������0ҋ`X�R�_4,-��m#L�ai�+�?���6�����RS~Az1�0��i�
�x7���,4\5�!��4�9\i+�{~�1��o��)�Ӭ��Z����wNu6�H�k�3p:�;z逭���]3ΧB)!t��,/&�J_�KG{̴y��m�h<�>%����$y��3���V�]%i��#t��n����V��J�7IZF (�� � r� 9@�ZT V�<��יZ�#^daǩ-y���20��F���יZ�#^daǩ-y���20��F�¦�T�#
��aSP�*j�MB0��F� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��6���9ClP��5�¦�T�#
��aSX�*k�Mb0��F5��P�#
�aCX�(k�b0��F5��P�#
�aCX�(k�b0��F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F;���aC�P�F;���aC�P�F8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x;���aC�P�F;���aC�P�F&���`�i�q4�8�lM6&�M������aC�P�F5�
m[k�/U�;��Ŏ��uɴb��1rm�z�h^���Íb0�Xyz�6�\�F.M�;���N�'�����������r��z�\�x�^�W/^+���׊�੬x*^�W/^+�o�I��$��m���x�k�[g�ơ�e�Fm�	Zǉ��yz�h^�W/^+���׊���r��z�D��k���b&��z�Az�A�x �<m�6�ǋǋg��]�u��]z��_����<X�<X�<X�<m�&�p�
�4�@ :�N�#:O����Ʊ�Ʊ�Ʊ�Ʊ�Ʊ�Ʊ�Ʊ��X�A�x�m�(�g��⩨x�j*���*�¹��t���$aw��d@�8�<�H��3����2�<�H��0����7�q��c���7�`����т��0SF
U���p�8t � ] .��A� �ŀ;�.��t�׷L�{,��h'L�rtχ'L�rtυ���X>���`�[zO���PzO���PzO���PzO���PzO���PzO���PzO���PzO���P,e��l�V��
���Z�X+S�%j���Po�֛V���a`�Lo���h~X>���j��F���j��F��Z�e�k�%="QS���aț���!�����r5��1���Љ�yǞ�I�]�
�zJ;��(� ��X�-�H�Φ�9m	�婵�鸛U��ګ��jGY�i�U}ze%xW�%x���8Ɲ���,g�"���D��U&X�c��Q�4�\9e�Q����B�8eӇ��[�F�_��Ŵ|߈X�����gN�1�#�>|ʯ���a�ر����?���c�y�?�i���q��݋,J���%��0i�|W�X��W��˧o�o��`����}z��-���zOM�#�u���(��;�/�4��ċ�Ų�?Ų_0A ��2�_F������?4!h.ߣ�9�G�j�1�j��+-Ĳ�ڙ��6��]:�������t�V�Ө�GL��ЊH�!������/'�h�- �bP��h@�>'�̭y����H�����H�+Q�����V����O09��#t��n����|:O�'I�D�>�'���@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9CP�j�mB�M�V��
�6�Z&�+Dڅh�P�j�mB�M�V��
�6�Z&�+Dڅh�P�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��i�Mz&�^���A�נ�k�q5�8��Mz&�^���A�נ�k�q5�8��Mz&�^���A�נ�k�q5�8�mP�F&х	�aBmP�F&х	�aC��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x;�N�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�S��T�x8�N7�SJ�*iQ�M*0��F4�¦�Tң
�TaS\P��5��p9C\P��5��p9C\P��5��p9Cl�hk��h�N�	�b���y�!�@���ƅ�1�z�h^���Íb0�X�8�#/Q��uK�uI�b��1s�����D�x"w<;���N�'s������D�x"k
�ǂ��੬x*k
�ǂ��੬x*k
�ǂ���r��z�\�x�M��&�j���V��q�xjZ�aơq�x%k'�������z�\�x�^�W/^+���׊�๬F"k�����ǋǋg������X�cl�cX뵎���^����z���5�6�g���ۮ��q���?5�N4��x �+U5�5�5�5�5�5�5�5������l�\�<U5MC�����@�J x�<N:H��;��<F5��C�ȁ�q�x�y�]'�;��.�т��8������7�`����т��0SF
o��M�)��:ekۦV��ekۦV��ekۦV�t��N�Z] .�C��2���+^�2��]|>���פ�[zKE���NzKD�uh�.��բp��PzO���PzO���PzO���PzO���PzO���PzO���PzO���PzO���P,e��l�V��
���Z�X+S�%j���Po�֙`�l�����X-���`�>V�Quh�V�Quh�tģwL�-zD���J*zD��L9tÑ7�9zC��NCF�r5��1�]�:g�y�<��H
$逮�����2��zJ:H9n
GN�N��o�ьއ-M�M�گN��^�R�1�"�~&���)+�~W������\iڑ�i��!�7���+��?�/F7�-�wU�m��~H�e�CL�#C���	�"X��l�q��7�,?�-��2-����7�w|ί#�g��L��w,E^ic���o�,E�)c��/�?�,x��~#�E����wſ5y��5���B����b�8��|?�o֤4˧�2�C����h|��Qƚk�/�U��<_0^3ТW�"D[�1n87"�?4'�o���ߦ99^��Uz�Jo鸚]9�Yt͡�N�h�u5�IGoC�4��u#��EЊH�!������/'H��y��o2��%:O�I�@�>eh�`�,�m��H�������V��J�7IZF�+H�%i��"t�N����|:O�'I�D�+D�eh�̭y��o2�M�V����7�Z& (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P (�� � r� 9@��@P�+Dڅh�P�j�mB�M�V��
�6�Z&�+Dڅh�P�j�mB�M�V��
�6�Z&�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�^���A�נ�k�q5�8��Mz&�^���A�נ�k�q5�8��Mz&�^���A�נ�k�q5�8��Mz&�F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F&х	�aBmP�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P�F;���aC�P��5��p9C\P��5��p9C\P��5��p9C\P��5��p9C\P��5��p9C\PX^�b�X�.�V�^�L�����i��9����Zez�2�.�.�.�.�V�k�5�痨ƅ�1�z�hM�&�
�oI�����Rm�6�T�x*M�&�
�oI������m�y6�<�x�M�O&�'�oɷ�����m�y6�<�x�w?����s����m�%ڇ��0��]�xm�'��V��y�x�k'�ǉ��y�x�k'�ǂ�s����z�D�x�M��M��M��w:��<Q6�M��X�A���?�^�ؽu�z�c�������������z�D�p��(˦��^(�U�z�D�#&��6�g���l�D�<Q6�M��sl�\�<U5�C�����@�8 x�y�^g��IZ�����ۤ�~m������	���d@� F#��`qO21��V�:@�%k����t��:@� pΐ8gH1`�X+A
�E��`�X� �ł��V��ekۦV�zO��u��.�]3���>���9�-����P_
��@]|(��L�l:e�a�-�h�t�FæZ62Ѱ閍�L�l:e�a�-�h�t�FæZ62Ѱ閍�u�.���`]|6�������i��kL�|&����L,����]Z5EգT]Z5]1(����1(���ޑ(�����QC���!������1�t�:�d���H�#oH"6�q�L��;��]�
�zJ;��(�'�����Ԥt�d��ӧ1��婵�鸛U��ڷ��wW�YX[��|�J�����p63RR�3�КA�1��"ǃ~0��i��r���
���n/��ſr87�o��x ����Ĉ�+ȯK2-���q^R��+�ߊ߈X�^r����~W�r��i��R��~W�r�꼪��0X��+����y[�E�lX����R�E����#~��i�o�y���1�"���^����/3q|��CM;����-�����]cNu+�"��I��r����-Š��O��'?�������r�M/H�,�f�w[Cj.�M{�Q�פ���0�^u��y���E$X��r�y������t�OW�h���BЀ@� t��n��m�Z�ςG��H�>	�1���Z��Aיh:�-^e�̴#y��o2Ѝ�"y�Ȟ`r'���"y�Ȟ`r'���"y�Ȟ`r'���"y�Ȟ`r'���m���`q6�M�m���`q6�M�V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5��&�ZD�+H��iX�"k�Mb��z&�^���A�נ�k�q5�8��Mz�#^�ר�5�0�z�#^�ר�5�0�6�"M��o$���6�"M��o$���܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0��F5��&�D�#��a\�"k��Mr0��F5��&�D�#��a\�"k��Mr0��F5��&�D�#����h�|y�`���@9{w<K�Rm����|#�τu�cX��V�k��h���l�J��k�5�Ë�cB���z�h^��Q�ׂU�1�z�J�F4/^	W��ׂU��*���z�J�x%^��^	W��������m�y6�<�x�^��^	W���Ļl�.�<�����C��l�8�<N5��c��X�<�<O5��c��X�<�<O;�+��K׊$������s���[���๶x�m�(���c����X�A6�A6�A6�A6�Az�D�x�k�ǂ�s��3�+��8�x�q�k׊&��6�A�x.j�����๨x.j������x@�J x�<N'g�Ǚ�1�x�t�"�dc�V�o��21��x������H3̌~y���21����t��7�h�� �ՠ��V�o���Z��@7�h�� .�E����}_���]V����1uZ����I�	�>]:���-�2���-ޒ�mӒ��9)=�-�h�t�FæZ62Ѧ閍7�Ji�"SM��oH��zD���%4ޑ)��M7�Ji�"SM��oH��zD���%4ޑ)��M7L�l:e�a�-n�h�,�2�h�,����V������Z����uh�V�WLJ7tģwLJ7tģw�90zC�N9(t㒇L9tÑ7�9zC��t�:�(�LC$zA��zA��z@Q'Lw�`+��(�'N���)�;pS�vвt�d��BiӘ���n&�zu���c����;��S|����
�D��<�C��b�m*Qm|����O�
�/F7�k���&�w����!`?�2���b-�ԅ�Wס�9c�3�%z���3�,|���_��i�����*�_�;W���c���Ƙ,~K��X�K��,~%���?%�U�?U濻?K�:,r�*�������?�?�h����W��˧~4�P�1�#\X��ŰM���W�]!���٩���n�iHo�֏�
�Ɯ �W��j��IJ����[��f�zf����&?���Lq�r�JΝ���3h;����N�k�nG����0�^u��y���E$X������)~����)��D�bP��Jy�C���@��D��@�-�%����$y���2�u�Z��Aיh:�-^e�̴#y��o2Ѝ�V��J�7IZF�+H�%i��#t��n����"y�Ȟ`r'���"y�Ȟ`r'���m���`q6�M�m���`q6�M�V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1���V�5��&�ZD�+H��iX�"k�Mb��z&�^���A�נ�k�q5�8��Mz�#^�ר�5�0�z�#^�ר�5�0�z�#^�ר�5�0�z�#^�ר�5�0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0�܌"w#���'r0��F5��&�D�#��a\�"k��Mr0��F5��&�D�#��a\�"k��Mr0��F5��&�D�#�� I�pMB��@9[,+m�
���.m@���Z=���A(�h�Z
M����:�Z1�V�k��h������Ze6�2�8�FM��M����&цS`�h�)�a��e�Fk�Z�a��e�Fk�Z�a���*m�6�J�x^�5��-b0�l]�x�j�q1@�G#ڇ����q��k�Z��V����x�k'�ǉ��y6�T�x�w<W;�+�o�I��$��m���x*k
���������m���Z&�։6�D��^�W/^+���c�SX�T�<&��dcCPyz�\��^�W5�K׊!1P��@�h<���@�J x%<N<��3�c���<E:ON��S��~j����x<_�$`u�����g�gI�F t���;�{o��e��Zo�@M��������������������ȰZ9G"�h�X-���`�[tχ'N�vt�Gg��[zKE���[t��NJOt���Ji�"SM��/H��zD���%6E�Sd]%6^�)��M��Jl�"Se��/H��zD���%6^�)��M��Jl�"Se��/H��zD���%6]8���-�N9n�q�u��1)1��1)0]%���uh�V�WL�-t�BפJ*zD���90zC�N9(t㒇LC(zA7�C"zD2'�9t�4k�!�:b#��� �����w��Ө�n�
�t�W{�Q�:����ۂ�9:�.��,���t�3z�3��n&�zu����;����4�񪾎$��W�"�|恧|�b���Q�No��V7��$��A��q���^��^f�4Ⱥ7�_8���,A^��~4Ӥ���(�,pX����ŏ�W�X��;~Q�7�`i����[�64��e���F�,r4�~R��Ƙ,li���X��)c��e���W������rǛ�K�c�̍��������~Gs~ Ӆ_3���-�r��2���"����hy�yŲ%7��?�F�W�ɤW�ҰW�q�|���B�]�C���ɏ��'+�j�����jf'L����jt͡�t����ۃz��tӦ�ŃΧo��`Cp7�������.��9w�C�'Hr$�D�!ȑ`J,	BM��@��D��@�-�%�ۤ�y���2�u�Z��Aיh:�-^e�̴#o����o����o����o����y�Ȟ`r'���"y�Ȟ`r'���"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"j�MB���V�5
�&�ZD�+H��iP�"m�m����|�ς6��F�>�g�l�#m�m����|�ς6��F�>�g�l�#m����Z�m����Z�m����Z�m����Z�m����Z�m����Z�m����Z�m����Z�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�^�ר�5�0�z�#^�ר�5�0�z�#M������`�i�r4�9l�6F�#M������`�i�r4�9l�6F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#k��Mr0��F5��&�D�#��a\�"k��Mr0��F5��'N�ޒ��t�S�Hr�m�M����!���@@Csj/�@��������P��(Rmh��>�g�;l�Gm��b�cX��+F/A˯A˯A˯A˯A˯A˯A˯A˯A˶���`r�9v��l]�.��m�˦�)So�ׁ����X�2��j��h���]�x#�`qO08�1�xm�'g����q�x�m�'g�V����x%m�	W�ƅ�1�6�T�x*^�W/^+���׊����<5MC�Sl�\�?�6���c�m��z�\�x�^�W5�Mc�SX�T�#ǂ��੬x*k
�dcCX�T�<5�B�@��@�h<���@�J x�y�#g��I�)�x�t�"���3xo� �C�P����<<� �3�1`���ƒ��t��$`������h"�Z�V�,����`J},�ł�ذZ;Gb�h�X-���`�r,�E��ȰZ9G"��X>ޒ�l9%9�rRs�%':rRpr9OG*��Aӎ[.�r�t���]8���-�L9n�a�uӎ[��r�t���]8���-�N9n�q�uӎ[��r�t���]8���-�N9n�q�t9!�$4�䆘������Oސ���O��Q��]1(���ޑ(�����(����9�Ӑ�]8�9!�� ���yȝ8D�ӄH�9��h�LC$zA��zA�N�:g�yӁ]�IG_�%~�ۃ�9:��$���b��B�91����o�9�އ-L�����^�m��:����4�q�����H�U�Hi��c�����Q�%�i��V>`*�,HQ�4Ӹ"��Xu?��m�]8�-����u�8Ӈ��%6��^G��0i�xo�|����b�e�?��8�¼�L?�W�4����W�i�y[�0�+~UyU�W�^UyU�a^Q��6ߔi����7�`����别�o�p���*��������~Gs�����X[z4<.�6�1�����?�ҁE�!�d<��b��B��m)|��>5�u~vW��=^��%z?���'?����ڙ��ŗL�6�H�k�;po^���t�V�]�K�N.�RE����/&�9y5�`C_��!����9G e�(H�����J o��J o�H��t�H�H��t�H�H��t�H�H�:��K�4�Z#K�4�Z#K�4�Z#K�4�Z#]%i��#t��n����V��J�7IZF�+HڅiP�"j�MB���V�5
�&�ZD�+H��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>��1��@�#>�g�l�#m�m����|�ς6��F�>�g�l�#m�m����|�ς6��F�>�ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�[ej5�V�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�Z�qְu�k�S`�i�r4�9l�6F�#M������`�i�r4�9l�6F�#M������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q�������a\�"k��Mr0��F5��&�D�#��a\�"k��Mr0��u��	Mפ�]2�`��n�w$ڵl@CPSڀ��lvk`�����(��)zJ�-5��C�3l�~m��Ͳ�����k�5���qM`8��SX)���m�˶���`r�9v��l]�.��M�R��)W��b0�l]�V�>��v��1�x����v�SP)�F#���c�b��qz�8�x^�/^��ׂU��+X�8�#/^	W��ׂT���X�<�<O6����+P�<�<O5ͳ����6������z�h^��ǉ��y�x�m�	[g�V�qz�h^��g�Q 9��q�x%j�<���20�̌<�#<�Ï20���2�<�OwI�)�x�7��f����/e��`��<7�c�F>�������я����߯;M��[�1���K wb�ذvU�b���]%9���1t��.����S��JsIKb�)l]%-����uh�.��բp��NV����9Ӓ��9)89��#���r���m��Cl?�aӎ[.�r�t���]1)1��1)1���`rCLHi��09!�$4�䆘���`rCLHi��09!�$4�䆘���D��O�8D�ӄO�9�Ӑϝ9�Ӑ��1(����1(��L�(�ӎJ1���9�9�= �����w��Ӽ�N�"F�㮘"�t�k��� �����w��ӄG�3�<�������;py'S�ӝN �$��hR?�ФLf�91��Nc7��SkC���F9�^��zc�E��KW��D4��<i�⸶�
a�jF�m-E�&�סX�����!G��N���M�ho���v�.�Z|4����&��[E����6Ŏ��/���0�9��~�?�W����eyU�W�^s�
�U�?��5^s�
�U�?��4i�y[�0�+~Q��W�^UyU�W��+�a���,t�5������7�o�,D�����7�k��<��^�ثѠ��u鿲��M/Lal��Qm������,P�A�[JE_�+�1n�������?����LF99ӝe0帕���bt͠��Cj􎦽ӷ�ӷ��[�u�Y �I��`Ct7A`y7���!�������`m��.�@����9,	BE��x��7�Q%:D�k�JF�D�k�JF�D�k�JF�D�k�JF�D�k�JF�D�k�JF�D�k�JF�D�k�JF�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�A֡h:�-Z���P�j��B�u�Z�A֡h:�-Z���P�j��B�u�Z��F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C���|5��kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F�U���h��Z:�V��U���h��Z:�V�����`�i�r4�9l�6F�#M������`�i�r4�9l�6F�#M������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q������`�n0r79���F�#q�����&�D�#��a\�"k��Mr0��F5��&�D�#��a1��'a��i`����L��
| !�:A��"� !�5�ֱh���/V�����P�{j g����V�m������l��>�ehf����+C5����Z�V�6���`r�9v��l]�.��^��o�.7���ĻX��#�
����|k(��SP)���j�6��v��1z�8�x^�/^��ׁ������q�.��k�Z�a������q�x�m�'g����q��k�Z��U��l�<�u�^���������x�k�Zǉ���q�x�y��/]g�n���e�V���ڇ��0�P�2�#5-C��P�2�<��C�`��(@�~y��g�g����<:O N���|9G!uZ� F?���N����*����� �n��ذso�1uZ���b�)l]%9����t��.����RغJ[IKb�)l]%-��D�uh�.��բp��NV��Hr��*��A�T����m�zCn�$6��]8���-�N9n�bRc�%&:bRc�%&$4�䆘���`rCLHi��09!�$4�䆘���`rCLHi��09!�?������p�����r�!�:r��!��bQ��%�!Ƀ��:q�C��:bC�!�!��"T�"n��"t�9�yȃ��t9y�]0E�(פzA��t�9��:g�x9Q�<�;py'S�9m	'�c)��hR?�ФLf����1����M���ڿ�ԯLrʽ1�#H~%�����~O,a��4��iڑ�[_$�����u>`*�,HQ�4Ӹ"��l��7�i��_��B���+�|����~Fر��W���-�~j�>dW������m�_�+�4��cL7�,a�)c���K��W��ʼ�M��m�*�Ѧƛm����+�ߕ���-�U�9`��~V�V�/���Ų�ݿ r��i���8��W���*�h,x]zo����Mchy�y�����0^8uD��2�_[J��G��|���zf��?���LF99ӝe0帕���bt͠��Cj􎦼9:����7�IGM�:Ȱ�ЊH]����!� �Ȱ����!�������`n���G b��]���"�r<XG��(��Z�D�k�JF�D�k�JF�D�k�JF�D�k�7��#�7��#�7��#�7�� ��F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b���F |�b�P�j��B�u�Z�A֡h:�-Z���P�j��B�u�Z�A֡h:�-Z���P�$j�C���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#X�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���kX�F���j�Z:�V��U���h��Z:�V��U���h�l�6F�#M������`�i�r4�9l�6F�#M������`�i�`���F�#q������`�n0r79���F�#q������`�n0r79���F�#q�\`�n4`��ƌq���у�0r70u�F�F����h��9���F҃����m(9JF�#q�����&�D�#���1�0�|�#k�ms��|�##���1�0��;!�Ƶ+p+��]dMb��Z��r��[ejx�9PTv�~�����7!�ͨV�7��sX�vk���ó!�<�&� ��\@�}k�mC�X�{m��k���Z��>�e����Gy����;l�Gm���`8��;�l��+C6��`p��3l�    V���@8��SP)�F#���v��1�xkǀƱ�1�xkǀ����#�db;l�Gm���1�F#���v���#�db;X��<5���ĺ��]z�8�x^�/^��ׁ��ĺ��]z�.�<5��c�cl�Gm����Sl��<6�MC�3P��<��`��@� F#<��0;����+]�����V�:Hŷ�Z���ӛ��9�-��@]|(7��p��Po�D�u��։���@]Z'��t��.���Rۦ%'�bR{�%'�!ʃ�%'�!ʃ��=!ʃ�!�9���m�NCl:q�e��!���-���t�:c���p�����p�����p�����p�����p���!�:r�!�:r�!�:r�!�:r�rj�!�rj�!�rj�!�rj�!�rj�w����v��yڮ��j�w����&�"`��&�"`��&�"`��e���Z��e���Z��Ò�rCHboH�D�dOHr:�#����t�4k��� ���!�:p���:g�x9Q��IG_�v��t����Χ r�OI�,]9��MM4��f�9jmk�n&��u���Yo��įG����HZ!(�ho�:�,KБ�Mj-�e��-������-���n2��a��ˤc�2������ԋW��b"�,o�oȽ~�#�,v߄[K?�o���c��E�[��l4¼��g��L+�a����?�ߔi�y[���c���,r�¼��[��o�4ڼ�M��l4��g����7�,pX�����W�������
�#|߭I�#���t�w�é�#\9x(-��ſ7�&-�B�^&�_[J��G��ʾ�u0r8���pBW��091ơ�q+=#���A��6���M{�mGLu7���oE��,u �X��U�y���p7A`Ct7C�������k����,k��9w��!��C�'Hr$�D�bP��J y�D1(��%<Ģ��@��e��̴y���2�u�Z��Aיh:�-^e��̴y���2�u�Z��Aיh:�-^e��̴y���2�u�Z��Aיh:�-^e��̴y���2�u�Z��Aיh:�-Z��#P�$j�C���|5�F��H�>	��#P�$j�C���|5�F��H�>	A��l@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-ڇ�#P�$j�C���|5�F��H�>	e�#l�$m����Б�Z6�BF�hH�-	e�#l�$m����Б�Z6�BF�hH�-	����:5z�^��W����:5z�^��W����:5z�^��W����:5z�^��W����uz�^�GW����uz�^��\h��p:5�x�es���Z5�A'0u�x�eGYBmZH������p:56�$q�\h��p:5��w�Z���&u�4��(8�J�$iA�ZTa#J:ң	Pq֕H҃����F�u�F4��*0��q�����c��J�#iV����uƌw<�h�֕�Dx��*���V�����L(�$
#	��@�0��6��#�����xת1��AWYṢ�����W����N���r�y���js��U�h>Tv�`l7��A�Z-�Aݗ���Rq`l5��6����>�Š%���z�{^� 5���)��Z#�AMB�SX�~k���p`8�X�Fk��`p�80 �0�0�Z� V�5 ⚀qM@8����#�ǀƱ�1�xkǀƱ�1�xkg����)�x
m��g����)�x
m��g����)�x
m��Ǌ;X�G^��/_�ǀƱe�xkǀƱ�1�xkǊ;X�Gk(��Sl��<5 �C�3X�{kmc��x=���M�0P������M�0l���� �@;�Z� V��� �mB1ɨF9��ejsZ(��Z(7���Z(7���Z(7���Z(7�����NV����9���1)=��ސ�A�T��A�T��AӐ����t�6�ri�!��!�="c�!�="c���p��r�/9���p�����p�����p�����p���!�:r�!�:r�!�:r�!�:r�rj�!�rj�!�rj�!�rj�!��yڮ��j�w����v��yڮ��j�p����/9hr�/9hr�!��"T�J���S��?����?�����p��!�]9�I��#��� �ۧ�:p��r�= (�r��ޒ��t����ۃ�ӝN �$�9��t�2�����1��婵�鸛_��wW�9e�G���N�~�/L�-��ib���c>M�����Nq+��-����7�&ߐB�o��_�M�J�<�X�.�Zo�ߣ��*�ı�����&��+�.��e^�_�>f`���q���,tߕ����a����W�����o�4¼��F�`����+�`i��ƛli�y��K��l�(��Ƙ,v��^ab/�7�?�߯���B�h��x2߭I�#���t�w��f�ߑ��$|�o�<�|�Ux-�B�_ �⾶���b�>Sp��� �8!+�����P帚^��YzM���Cj􎦽�6���:��u�&���,u �X��U�y���p7A`Ct7C�������/"���,k��9w��˽����!ȓ�9t�"O1(y�%<Ģ��@��bQ�J y�D�)����)����)����)���2�u�Z��Aיh:�-^e��̴y���2�u�Z��Aיh:�-^e��̴y���2�u�Z��Aיh:�-^e��̴y���C���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j��؁h6 Z��b�؁h6 Z��b�؁h6 Z��b�؁h6 Z��b�؁h6 Z��b�؁h6 Z��mC���|5�F��H�>	��#P�$j��Б�Z6�BF�hH�-	e�#l�$m����Б�Z6�BF�hH�-	e�#l�$m����tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�h��Z:�V��U���h��Z:�F�Aѭs��6�$w�G��6��:�V�8դ�56�$k�m+ĉ��q�B������x���m+ĉ�x�8у��tjmZH�|�_m*0��F4��F�Hң	Ta#J�$iQ��*0��F4��F�Hң	Ta#J�$iA�Z�a\P>|�Dm*Ѝ�Z#]����0u��6ġ��H/F#Cβ ���^�D���A9 �6!F��V��ڔN�rp��词�Ig���7p�]:��;q$t�1�7y�)�1)��|=����GOt���.�鎐� Z6ej{l��+S�jմ�����{w- ;�����B��P�{k�mb��z�{^�ת���8%��z�}m��[`w֡Z������2�P� �+C6��Ͳ�3X���5����`��0R�)z��F
^�/Q����K�`����z�~^�������z�~^�����F^������Rm�)6��x#���c�cX��<5��c�cX�Gk(�c��x��������<5 �C�3P��<�ǃ�l��#6��M@;�P������M@;�P������k��Z� V��� �mB1ɨF95�! :ۤ�Oo�E���,	M����,	M����,	M����,	M�uh��I��I�Hr��*Hr��*Hr��*���t�6�ri�!�ri�!��!�="c���p�����/9�r�/9�r�/9�r�/9�r�/9�r�/9�rj�! �"`�L���r0B&�D�9�! �"`�L���r0B&�D�Ӽ�WN�];��t�;UӄL8D�ӄL8D�9y�C���9�!��"T�J���Pr*A'�"A'�"t�7N#t�4k�!�^�Dm�F�;�@��rN^q ��z@Q �G_�%~�ۃ�9:��hI-�$��e#�1����o_ьއ-M�M�������1�-�?����bGhr����_���|WѠ�X�1�i��"�|�-��
��W����%�%?��n��ı�L2�C��U�&-�������?�W�]n4ʼ8|����f�Uy��F�o�W�ߕ^V���[��W�i�y_�o�4���U�0�¼Ѧ�W�4��
�K�64ڼ����W�4��g����7�,v-�b[��o��A�����>,E^�L������M�����l���e�+[�8_0^3ТW��j��IJߣ��[��a�����pBt�I^�İ���-���b˦:�N��6�H�k�1�޺c��[�h�Qԅ���@�t
�o�;�������,n����o㗓�����X��~��.��9w���9t�"N��I�%<ġ瘔@��bQ�J y�D1(��Z�KA�Ih6�-�%�ۤ�t��n��m�|<ςG��H�>	g�#��$y��3���|<ςG��H�>	g�#��$y��3���|<ςG��H�>	g�#��$y��3���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C��@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-�A��m�|5�F��H�>	��#P�$j�C���Z6�BF�hH�-	e�#l�$m����Б�Z6�BF�hH�-	e�#l�$m����Бz�^��W����:5z�^��W����:5z�^��W����:5z�^��W����:5z�^�GW����uz�^�G]���p:5�x�/_k���\�#�ȇ�kJ�$
<GSj�p8۸m6� i^#��\�F�n�ڴ��6�F5�k\�F���ׯ��h$ң	Ta#J�$iQ��*0��F4��F�Hң	Ta#J�$iQ��*0��F4��G0u�x��х�+�|�q���kB4���>��tj��6�Z�Q�b�YP��P�F�ħ�J�$
��A� ��T�I'/��K��R�6S#���%�Sh�B�r�p t͠�]mb��Z�ӗ��Kգ�P9O, ����@J?k�����/U���Òmh	6J{M�_��@�`�٬%9/V�n壚mZ�V��ծi�k�X�sk�B�٨V� �%h'IZ	�|=��C�l��+C6���`;�X���/Q����K�`��0R�)z��F
^�5���b03X��#5���b03X��#5���b03X��x?/^ɷ����Rm�)�x
m���1�F#���v���<6�M��Sl��<5 �C�0� @�  F m���d`&�	�}j�D
�a��@�vj�Z�w���@�v+]�gÛ��sy��M�h��>�ejs̭Ny��Γ�=��S`]����L]����L]����L]����M�-����*Hr��*���t�6ç!�9���m��"�B-0�"�O;e�<�N�:p�����p��r�/9���_�����W�j��+U�Z��
�@V���_����sw�󖿧���<���-O9k�y�_��Z��r��󖿧���<���-O9k�y�_��Z��r��
n�MÐ)�r7^r���-^r���-@R��*O9C�y���P��r���?���^��j��#W�9�y�×�t9y�C�� r$t�9�y�;�@�G���I�@��Ө�oIG_�v��t����N��$�ь�t�2�9jk'�c7���oC��ֿ��mGY�^����J�~17�LB�1�E&��CH>4+�inK�H�0u��A\ߛ��,H��JJq6����7�^��o�ߣ��N,A�����e���U�2������a�^{~Q��K��64��cM�6ߕ^k~UyK�6��~Q���o�ߔi�y[���c��Ѧ���`��~V�V���߫�W�X�c�l������t��`-����W�`�*���dt��~�?���6��n2bG���]b�_8M ��D��v���������������ɡɎ5t�L��b˦:�B��mt���鎦��M��E���o�U��X�:��������!����^M�r�o㗑`C_�5��������`n��I��:C�'��<���bQ�J y�D1(��%<ĢIh6�-�%�ۤ�t��n��m�Z�KA�Ih6�-�%�ۤ�t��n��m�Z�KA���H�>	g�#��$y��3���|<ςG��H�>	g�#��$y��3���|<ςF��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C���|5�A�l@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-�A��l@�-�A���H�>	��#P�$j�C���|5�F�hH�-	e�#l�$m����Б�Z6�BF�hH�-	e�#l�$m����Б�Z6�BE�:5z�^��W����:5z�^��W����:5z�^��W����:5z�^��W����uz�^�GW����uz�w�]�����Mz�m�C��th��Fx���У�u�x��ф����X�w����������]n	'I�y5�A&���?��&��:�<�*0��F4��F�Hң	Ta#J�$iQ��*0��F4��F�Hң	Ta#J�$q�Z�k�Z��5�A7(��J^�	j�A�L|�#iA�\o�k���M���`��6҃���B��A9!e+0���<�ܒw$�^��y��G'�����N��P��u~�W��5��m��5����=z�n��)j�jc����>m�Ѱ�-ڂS�P9}m�/k��%��9�JPq��kD���=��Nw>���&�Z��+\څk�P�v+]��N�����+^څk�P�{j�m�8�X��#5���b03X��#5���b03X��#5���b03X��#5���b03X��#6���`f��F^�������6���5���`;�X���5���b03X��#5���b03l�Fm����w֠��F;5�f�� s����ek�̭r���� �o2���V�:O��I��>�0E�.�[��)��֍6��i���`Jl����`Jl���`Jl���`Jl���`Jl����9i�����9i�be��/H"�zA���^�E��-פn�w�1Ӽ鎝�L@����9yϝ;��t�;T9�� Sp�
n��s��� Sp�
n�MÐ)�r7@����9���)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��?�)S��+�(�����(����ל�^��j��#W�9�Q�_Ҏ:�����F��*5�Q���O8�r@����$���n�Gt�8r���pz�v��t����N����hI?�N�5�r��O��o_ьއ-M�M�������1�-�?����b��	^��W�&��CH>4+�inE�,�o� �xF��y�ߌ(�q�Ciz��:G[~N-"ߢ�b��+�o�X�������.�^`�*�ߊ��i����o�4�c������li����6��~Q���a^j���7�W�����M�ʯ)c�y��?�6��i��+�X��9c��M�ۿ���J�+��M��b�K(-���MI�(����t�q��é���0�;���Ŋi5Fqq�f�C�3~��z���q)#�1���Nu��;S1:f�wt͡�N�k�nGLu7��pM
;|����X�:��y����p7���X���X��r�o㗓����!�������.��9w�D���9t�"N��I��:C�'Hr$�G�!��9t�#�1(��%<Ģ��@��bQ�J y�D�؁h6 Z��b�؁h6 Z��mC���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C�m�|�����6�>ڇ��P�jmC�m�|�����6�>ڇ��P�jb� �h@ Z�� �h@ Z�� �h@ Z�� �h@ Z�BЁ�Z5B�h@�-��P� j���m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�k�tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�h��Z:�V��U���tj��F��ѣ�����6�%���m*0��iQ���Q�:ң	ρ���I�k���%�-Ãkn	!��M���h��F/u�#��5ƌq�\h��0uƌq�\h��0uƌq�\h��0uƌq�\h��0u�x�8�N5iC\�iV�m*�ҫHPq��)~҃�^����51���u����h��:>V�G��iLy��"�����Pڣhڣ��S�)dy�niF�dp��D��qp��}$�"�F���H[���u;����.������bL@CPy�i�18@Csm�+m`尛��c�����w�	��zmh��-�gÓl�r>��1���|9�χ7��� |>5
׶�Z��+^�`p�8�l� ��m��6��`p�8�X��#5����x=����c��Fm���`pc��Fkk׃���z�~k���w���~kߚ�w��Fm��6��`p�0P������k���@� s����'�Z��+\�'��̭ry��O2���|-�O��I��։��h��Z���>t�4�tr�G-�tr�t�4�LCLG-�tr�G-�tr�G-�tr�G-�tr�t�6˦!�]1��-פn� �uӼ鎝�Lt�:c�y�;Θ��t��
~�O�Ҏ|���P�
n�MÐ)�r7J9��Q�Ҏ`�[�k�Q�Ҏ`��s���?���(��G0J9��Q��P�Tr�z��+��^��
�G(W�9B�Q��P�Tr�z��+��^��
�G(W�9B�Q��P�Tr�z��+��^��
�G(W�9B����(�����(��y����F�^r5z����W���TrEz��+��^���
@�@��GJ8�����(r���pz�-�����{�n ��t'S��6��1�����C���Z������1��婵�鸛_��wW�9e�G���CH?&+�~RW���4�8\[�r�Q�o�-E��$�W?�I���F�k�/�/[��/3qe�=1lU��-�ӄ�|�y��~G�w�Β��ǆ�~*��č0X�����������ߕ����a��y_�oʯ+��[��4�~UyF�W�ߕ�)c��������+�������𿻫�i���E}o�i�>g,KP-�ӈ_�+�A� r4+�.���ſ��7�>�`^-���
������8���ko��lW����U�=�% �~%������r��jf'L����m,���7���B�pM
;|���I�S�:���RM��p7���X���X��r�o㗓����!�������.��9w�D���9t�"N��I��:C�'Hr$�G�!��9t�#�1(��%<Ģ��@��bQ�J y�D�؁h6 Z��b�؁h6 Z��mC���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C�m�|�����6�>ڇ��P�jmC�m�|�����6�>ڇ��P�jb� �h@ Z�� �h@ Z�� �h@ Z�� �h@ Z�BЁ�Z5B�h@�-��P� j���m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�k�tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�tj��F�Aѫ�h��Z:�V��U���tj��F��ѭ+ĉ��q�H�q���I�!��kA!��ƭ k����q���(�8D��klCw�դp8�J�$<��5�w>�kA'0uƌq�\h��0uƌq�\h��0uƌq�\h��0uƌq�\h��0u�F�>�U��h�
+Fŏ ��I�CX���
0lB:Ҿ	d���y�6�V����ֹZ�+Q�rIdm��%E�3�w�s��đB%�VYw������|�=&�D�yX�����z����_�1#�
|���e��(� ��<�6�Cl��6Ⱥ9n�C�Ȁr�m�-����k	M6�r�m�J�)@@JNj�mB�m�Z-�E��h��-�e��̴[j��B�٨V�6�ﭰ;�X��#5��M�;�l�����ﭰ;�l������b0X��#Z�`&���#5��ֱ	�F>���Mb1�z�{^�/^i���m�� ��m��6��`p�8�	�Fm���d`&���F;5�a ;���@��+\څk���� |9O2�m�Z-��E���@�ry��o2�m�%':D��H������+UӼ�Θ��.�[��)�X�"��.�[�����i�����i�����i�����i��r�tÖ��!�="c���p�����p�����p��r�/9�r�?�+U�Z��
�@����Z���O�
T���J�G(W�9B�Q��P�Tr�z��+��^��
�G(W�9B�Q��G"o���Tr&�Qț�G"o���Tr&�Qȕ�M^�D��M^�D��M^�D��M^�DÕ�9Q��L9Q�ÕL9Q�ÕL9Q��Ҏ:��q������u�(��G@Tk��U�H�TrEz��+��^�H��9Q����(�O�G[��9nP�G_����M������9:����N�C�m�c)��SX�-Md���|��f����r�����M���;���ߣ��^��'��ɮ��_дLo��D���]_��i�e�c>Im��0W?��<|7�q���6͡�)`?2���l_4X�b������4�?�W��;|4��߫��ر��
�W��+�f�W��+�`i���W�^V���[�64��e���F�m����F�,|ߕ�[�O��;�[-�����v�n�����e��(y����zC��M�~i�je�w_0%0y�-���CNo�����ܫ���U�=�A'�8�������P帚]9�Yt͡�N�i`���ދ��4X(��`����
�t�u;���E$��wy���X�����/&�9y7��ɿ�^M�r�t�.�Hr�t�.����y�OW���t�`n��!��D07H���� ���y�D1(��%<Ģ��@��bQ�J y�D1(��%<Ģ��@��bQ�J j�C���|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$m�m��m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�j�BЁ�Z5B�h@�-��P� j�BЁ�Z5B�h@�-��P� j�BЁ�Z5B�h@�-��P� m�m��m�|�ρ���6�>�g��l�^�ׯ����mz�^�ׯ����mz�^�ׯ����mz�^�ׯ����mz�w�������n�q�p8۸m�6�w�������n�q�p8۸m�6�F�U���h��F��Ѯ�tk��F���A��x����b���e#PCy]c�5i ���
<GZ�q��H/u�"aG���Fx��#�*0��q�Hρ�s�yƌq�\h��0uƌq�\h��0uƌq�\h��0uƌq�\h�֔u�<�>�����H/V���#�7[�,�z��t禥7	�I��&�h6>V�ZPq��(6�F�քn7�5��$6���Hޒ-�íx�Ƽxcz6eb&��H���S_����'�.��ѱ�%FN(γ�_�A��X��SgSu�n֡Gl��*`��b���]0�����d@9l�m7���y�)�Rp����-څ��P�[j	�C�=�|(5�����+\څk�P�sm��[`wf���F>���M�;�l���6�ﭰ;�l���6���b1��F>���ֱ��#Z�c�X�}k��b1��F>��������	z��x���/m�0l� ��m��6��M�0l���� �B1٨F;�� �b w7�Z��+\��!��@�ry��o2�m�Z-�D��h��-�e�ۤJNt�IΑ)9��S��)���s�?G-����o�F�Z4��Ѧ�֍7LCLt�4�LCLt�4�LCLt�4�LCLt�4ǤCLzD4ǤCLt��N?t����>^s���>^s���>^s��j��+U�Z��G0^r��*@R��*W�9B�Q��P߭�M^��
�G(W�9B�Q��P�Tr�z��+��i71��Ɠp#M��i71��Ɠp#M���Tr&�Qț�G"o���Tr&�Qț�G"o���7'����p"M���7'����p"M���(��GJ8��Q�_Ҏ:��q��F��*5�[��~���nm����Go�y�7����Ҏ$�[�r���pz����M������^�N���t'S��6��m�c)��SX����?���?��F3z�6��7k�:����,���bW����L8��8pKW������I^�b�5#Z�6�)c��u>`�o�X�o���M���c�+��B�~}"X�R��i_�?���>d|��J����,|��i��g���+�n�¼���0X�+�L9m�)c��Ѧ��c����_�?�,r��^{�����o�p��~�~�#�|�X��[���l*߄[�_2:p��3�?�����8�qm���x�0�\X�B�i��⾶�(��z���Z	7��#�,9�j��)�-���ڙ��6��]:���p:�;z.��`��ł��7�*��y���"�o��y���p7A`Ct7C�������/&�9y7������!˽���bS��%=^bS��!��D07H����"�Ct�"N�DI�%<Ģ��@��bQ�J y�D1(��%<Ģ��@��bQ�J y�D1(��|5�F��H�>	��#P�$j�C���|5�F��H�>	��#P�$j�C���|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�m��m�Z5B�h@�-��P� j�BЁ�Z5B�h@�-��P� j�BЁ�Z5B�h@�-��P� j�BЁ�|�ρ���6�>�g��l�m�m��mz�^�ׯ����mz�^�ׯ����mz�^�ׯ����mz�^�ׯ����m�6�w�������n�q�p8۸m�6�w�������n�q�p8۸mz�^�G]���p:5��w�]���p:5�
<GE�&�HXJuz?� *H(�F���{��^�"q�H��7s�y�q�HTa#J�$k����q��l|�F�_�b�Y�:�F�у�4`�:�F�у�4`�:�F�у�4`�:�F�у�*0���k��mq(H(�+Ho�椼w�
����:E0+���A�D(��r��|#SkB7���|8�{���0�X�*A$T����4�БSZH��@��@��yH��%'�D<�.=)��Z��Չɶ�6���b4���1ț`���� V�$17�m�LC?t�-7Hr�t�j�E�X�e��P�vt�o2�m�|'���Ѱ��-a)���-C�=�Z-�������+S��k�X��+\�ejsl�rm���b�ͬ[k�k�c���x9��i���m��x9��i���m��x9��i���m��x9��i���m�����ﭰ;�l������Ͱ;�l��#Z�c�l�rm��M�1ɨ[j�ڀu��8@�Ny�	�3�=�|'�KEIh��-g�{��Pt����A������o��`9i�C�ˤJn�D���7��a`C?,g���!����t"|.�O�3��t�;U�<�W�7zA�>t�;UӼ�P�
n�MÐ)�r7J9��Q�Ҏ`�[�j�n������TߧQS~�7����pW�Q�:����D߭���[A~��6�mm�������h#o��F߭���[A~����:���$oӨ��N�F�:���$oӨ�i6����ƓhM�li6����ƓhF25^�Dj��#W�Q�:���pF����W���[�4i6����Ƒ�@4���u#��iDH� GQ �:���7�ho��4�g��m�����w�������{�:���<��py:v��t�����C��6��m����S��N��e r��O��oU�S:-M�M���S�:����;�&9�^�#W��ɭ�-�~B|��$����_��_�n-��xX�7S�����օ�q��^F�?�2�C����F,@i¯���?�i�,|�˧W�4ʼ?��[%���7�o�,|߅�ر�b�?�a�ر��
�?��8�¼�L?�`����y���3?��`X���L�����[��i��X��]�ؖ0����|��=!��1`8�4�56����-���X��u|$�F�p�@�_$��m��́ʿ	:p�.�'N?�]8�MW�9L9n&�N���H�5:s��zGS^��v���VM�
�t�u#���'�N��)&�I7�����w`Ct7A`Ct7��ɿ�^M�r�o㗓�������/&�9y7��ɿ������t�.�Hr�t�`n��!��D07H����B��<�D�!ȓ�J-���l�$-BЀ@� -BЀ@� jmC�m�|�����6�>ڇ��P�y�C�1(y�%<ġ瘔<���bP��Jm�m��m�|�ρ���6�>�g��l�j�BЁ�Z5B�h@�-��P� ����(x@J����(x@Jj�BЁ�Z5B�h@�-��P� m�Cͱ(y�%6ġ�ؔ<���bP�lJk�bЁ�Z5�B�h@�-šX� ^�ׯ����mz�^�ׯ����mz�M�Ij�Dڴ�6�$M�Ij�Dڴ�6�$w�������n�q�p8۸m�6�M�Hj�p8۸mƌ$q�	h�G0���w�]���p:5��w�Z�q��mƭ �Ȝ`��r0�F�*:�Z�h��\T�#�a u�?i^m+�l&�;��N�h�J�i^m+�m�x�����6Ҽ�Ta ��T!x����m(8��F>F���jl�@��&�D7�#\�F���r��|;��(8�Q<�����0�(��I&�^\��v�b���������C
���C�a���j#a@q�c���}w�W�[���-c���"�,J-�����P:�ףQQ���j�bGK��'��%	:+V��&.Ԡ�6�X��HZt+��[��%/^	�H
n逧ŀE��-�Ln� �L]�7�R�`JOo���Jl5��l9n�G-��(�zJ?k
C�=�|(5���Z��+S��t�m�V������Z��+S��t�mz�[^����%�1�z�r^����%�1�z�r^����%�1�z�r^����%�1�z�r^��`wf���}m�ݛ`wf�ٶvm�ݚ�c�l�rm��M�1ɨ[j�ڀu��8@�N+S�g�{��Oy�	��A�Z(:KEIh��-%��%6�)���M��r�,	M�H��t�M��9Lo����~X���`C?B'��D�]�:g���v��yگH
n���j�w����&��9y�C�)���?���J�Ҏ`�Tr�z�[��	���T߭�M�[���no�	�Ө�^�DJ��"o��F߭���[A~��6�mm�������h#o��F߭���[@�~�D��u7��HߧQ#~�D��u7��HߧQ �mcI��&�64�@��mcI��&�64�@�~����m���[�����HߧQ#~�D��u&�64�@��:���@4���u#��iDݴv�<߭�y�[@��1��H�z�s~-�e��m�z����/��h_�өЯN�@ru:�����C��6��mzc$�ь�F2�9jk 婬�ьޫ֦tZ�Z����9n&��u����wLs��F���[�Z&p��-��j��}��ԛ��-F�&��M�7��-�x;~F�"��l��t��Ǟ��,y^�ث�u�8����?�p@����n4ʼ?��`X��W���7⿺|���1��b��+�w,A^s��b�b�9���eyϙ��,v߄�K>eW����U�%zX����W�ac��>ezO�^F�?���6����+~m*бE�|$Ɯ �,P�H� G�j����C��JN�&�&8��e`帚];S;�#������M{���d���'I�R:O:��y���"�o��y���p7A`Ct7C�������/&�9y7��ɿ�^M�r�o㗓���~��k�Hr�t�.�H����"�Ct�`n��%:C�'Hr$��`n��I�%�C�l@� -BЀ@� -BЁ�|�����6�>ڇ��P�jmC�m�%<ġ瘔<���bP��Jy�C�1(y�|�ρ���6�>�g��l�m�m��m�Z5B�h@�-��P� j�BЀ@J����(x@J����(y�Z5B�h@�-��P� j�BЁ�%6ġ�ؔ<���bP�lJm�Cͱ(y�Z5�B�h@�-šX� k�bЁz�^�ׯ����mz�^�ׯ����m6�$M�Ij�Dڴ�6�$M�Ij�Dڴ��6�w�������n�q�p8۸m6� M�H��n�q�0�ƌ$q�	h�G0uƌq�\h��0uƌiQ��*0�B�#$�`��գ�^�F���%��~/�C��4��^�#M� ׫G���:�Z=E�1�Đ|�$<I�A�Đ|�$<I�A��B�#k�����h�����Ta#J�$�ȅ�0��t(:ң	��k\6>jt��</x�"aW��A��|�Sjap�V׭M���N�@פ7{����8�D`ی��L`� g�_�n��§-�
�B����*�J)"�)�I	��(A�ao����$
�ѨܜA	M�*���D��3��Z6�Q�1ޣHq_�f�D�r��>t�M�tr�zO:b�n�I�5E�ʁ`CP,-1 ��[��Q���|�O�g�M�Z6g�M�|(5����Z��P^�S��ka�|(/A�����1=6��F'��ӝ�ŷr1m܌[w#��ŷr1m܌[w#��ŷr1m܌[w#��ŷr1m܌[w�/Aݗ����we�1�z�r^����%�1�z�r^�רŶ�9�Nm���=�V����ej�̭Py�����>���֍7I��o�F�Z4��ѦX�%�)�X�%�)���)���|��Gŀ�XZ���]!���3qt�n�&�"`�&I�-zO9k�y�^��Z��rפ�'��ӁJ�8�ӁJ��L9Q��L9Q��p"M�M�7%zu+Ө�^�Dj��#W�Q~����m���F���F24i�Ѥc#F���F24i�Ѥc#F���F24i�Ѥ�ƓhM�li6����ƓhM�li6��ncs�[���� �1 �1���@-�bz���hW��m^���z���hW�Q�:���7�ho��߭��[@~��6�m m�� �����hF3�i�Q�c=E�Sw�錿o�~�[B�^����:�
��t'S�9:����N��m���8錒F2�^�5�r��A�SY?��W�L��6��7hr�MO��;������w�?Ð�j�E�X�W�%}|��}	��.)���7%�Z�8M X������ň����A�����0������̯I��o��|`X�����~������.�^c�G�n4ʼ;,E�2��7�o�|�����~#�E�3��ߊ��i��B�>`��~�n߁�7�?��+�,J�[mb��1�E��#��2��M�0���4�n�q����U����AX4�4�Ӆ����T��87/�?'�p�.�'N8����5Lq��:�Ν�����jt͡�zGS^雁ѿ�VM�
�o�U���'�N�<�v�I7��I�������!����^M�r�o㗓�������/&�9y7��ɿ�^M�r�o㗓�9w�C�{�9w�C�{�Ct�`n��!��Ñ'H����"�Cy�"BP�P� j�BЁ�Z5B�h@�-��P� m�m��m�|�ρ���6�>�g��l�j�BЁ�Z5B�h@�-��P� m��Ͳ�y�V�6����Z<�+G�eh�l�jMC�I�|	5�&��$�>����P�jMC�I�|	5�&��$�>����P�jMC�I�|	5�&��$�>����P�k�Mb�I�Z	5�A&�h$�-�Š�X�k�Mb�I�Z	5�A&�h$�-�Š�X�w>�ρ�s�y��w>�ρ�s�y��q�Hj���ƭ q�Hj���ƭ iQ��*0��F4��F�Hң	Ta#J�$q�Hj��m�iQ��*0��F4��F��F�<��\�#<��4|�F���{��<�#�G��@҃�8� b�X�1|P�Z=G���0��#d�x1|P/�E��h����Ѣ��4^�F����{�,u��A�Pq�h<҃����6w�� n1�l��wޮ7���@!x�c�7��(� w-�ǝ���� ��H��0����cL:�w��N1�4*�?m���9��#
��7ش�>l�n�@~�3�/ڷ��$aI���$[t^F�k�/�X�*�
�"��N֣f!�D�D��5)A���^��f*�o��H]n+��c������D�"T�!��w���7��Cl��6�!�D��l9n�IG��Q���~�-��e�|4�g�M�|4��ka�V��ka�V��ka�V����u�1=6�OM����r1m܌[w#��ŷr1m܌[w#��ŷr1m܌[w#��ŷr1m܌[w#��u��Z������m`:�X������m`:sX���6����Z��+SڇP�Py��2�A�V�:O�ä�l:O��Z4��Ѧ�֍6��i���`Jl��Ⱥ9n����9L,-R�r�,-Qt�n.�������:`����:`���y�^��Z��r�N*t�R�N*t�R�N(t�R��GTq0�GM���7'����p"W�Q�:������ho��:߭�u�[@�~��Ѥc#F���F24[�2An���S$|��6���m�[�����n#o��F�5���kq|֦<��Ly�Z���1��jcϚ�ǟ5��>kS|֦<��Ly�Z���1��jcϚ�ǟ5��>kSo���Lb�1��� o���Lb�m������$4�a!�c=F���F3�i�Q�c=F���F3�i�Q�c=E�Sw�v��|��MM�4��ɿLg�~��&�m�m���8�hI?�ВM���Ld��1�J��I+֦�W�Mb�5�r��O��oU�S:-M�M���S�:����;�&9���7N8����&� �����]_����e}Ŋ�,�,�kЬ,aL[_ǋ~bib\o8�Ma��Ѐ�W�]G��H-���,`�~!bZ��CM5��3���zE��2����+�c��*�1�	b��o�X���W���%y��w�M��ey��&Ű����x2-���и��]zo�F;��a�ߍ�Cx|��{�_�5|	���,�+��-ƅ�~�sc��OHq:qĤ��`rc�]9�V[���53��1�B��mt���.������d���'I�R:O:��y���"�o��y���p7A`Ct7C�������/&�9y7��ɿ�^M�r�o㗓�������/'Hr�t�.�Hr�t�.�H����"�Ct�`n���^��"�o���C����h@�-��P� j�BЁ�Z5B��6�>�g��l�m�m��m�|�ρ��h@�-��P� j�BЁ�Z5B�Z<�+G�eh�l�m��Ͳ�y�V�6����$�>����P�jMC�I�|	5�&��$�>����P�jMC�I�|	5�&��$�>����P�jMC�I�|	5�&�h$�-�Š�X�k�Mb�I�Z	5�A%��yz�^�������yz�^�����s�y��w>�ρ�s�y��w>�ρ���ƭ q�Hj���ƭ q�Hj��Hң	Ta#J�$iQ��*0��F4��G��ƭ k����q��Hң	Ta#J�$i^#�+ĉ�x�4� ��t(�
<GB�֕�6!u��^$��a ��Hp���$o�L�B�$iAǅ��hy�Fp��c��a ��:/�E��h����Ѣ��4^�F����{�,x�E�@�9 �6,x�C���c�!F��.�p���%=Z�J�+G����0x(�z��'IGp5 W@A�@���'�@��0���&�p5�;�z�͒�����:H(9p���6;�4C��ۨ7bG�y��oy�����oy^F�j������Ĉ�Bu9U���k��MiT�:��;)�ƨ�HzvX�C�'�9(A��iG n�Sp#���k������l�i���"���mט��m�-��)��Z&&։��(��Z&5Dơh��>����>�b���>�b���+[-b���i�A�k�v�m��F'�щ�bzm��F'�щ�bzm��F'�щ�bzm��F'�щ�bzl9�[k���u��m�NkӚ�t�9�V������A�Pj���Z�>b�M�V��k`@�i�7�h�y����h�y���H��t�M�H��o���9L,g���!�����C0Hf���K]0D��K^��T��r���='��ӁJ8�9Q�ÕL9Q�ÕL9Q���p"M���7%zu�Ө�^�Dm��[����ho��:4�dh�1��ݩ�v�H4�@ط1���@-�b�jcϚ�ǟ5��+�qW��$���I_[����%}n"J��D����+�qW֦��L_Z���05}j`j���������SW֦��L_Z���05}j`j���������S�L[�01n��ŻS�L[�01n��ŻS�M�-ڛ�[�7x�jn�nc/Ź���2�[���n���ݩ�ŻSw�kq_�&��MM�-ۋ�[�@�jn����
��I+�$�Le:�1����S��N�Ld��1�J��I7�SS�֦�W�Mb���|���|��f�^�3�r�����M��q5?�������rc�Ñ����Hr[�_����+�|W�������^J��_%�ӇTE��/�F�,`���1��.�(�M�qi��ϙ]:�,y^��|>g�c�w������>goƽ~�������w�]3��y���y���y�����ƚj3�e�X�cŰ,P���}7�W�Ac�I_���o��P�N��~F��-�
0[C�|+4,�>j��|֤ۋq��J���À���OH~&:a���β��:�.����;S;�s��t���.��躣���
�o�U���'�H�<�wI�S���I��RM��p7���X���X��r�o㗓��aˡ��aˡ��b��!��b��!��7x������@Cw�n�� !��"�Co���[�E������(y�Z5B�h@�-��P� j�BЁ�|�ρ���6�>�g��l�m�m��m�Z5B�h@�-��P� j�BЁz�^�������yz�^�������y�Z	5�A&�h$�-�Š�X�k�Mb�I�Z	5�A&�h$�-�Š�X�k�Mb�I�Z	5�A&�h$�-�Š�X�k�Mb�I�Z	5�A&�h$�-�Š�X�k�Mb�Iz�^�������yz�^�������y��w>�ρ�s�y��w>�ρ�s�yƭ q�Hj���ƭ q�Hj����x�����6Ҽ�W��J�i^m+�m�<�k��r0��x�����6ң	W��J�
<GB�У�t(�
<GB�ֹZ$!x��$b��4B�do�u�V������X�Q�6҃�����5�I�^$���4^�F����{�/�E��h����Ѣ��ر�@/F�#`��AxD#I��#�����$8GA����H!k�K��EN�!�������R�X9X��b���S��,�
|)��JP/����>|�h(CY��{i��F'ӡ�M���a�����D��S����j��Z��z���w�0���9�T�ENP��M����I&N��Q��!�E��jImGm�6i�Z�O8\��#^�JwLc�����zF0��:���)��Qڮ�
|.���E0@?ji�@��@J?����(��Z&5D����m�����m�ֱZ�k���Z�^��נ�5�;M6�OM��h���1=6�OM��h���1=6�OM��h���1=6�OM��h���1=�V������Z��+S�ej{l�Om���=�V����Z�j��� |4������>b�L@�i��F�̴l��FˤJn�D���7��c�3���~X��Љ�>Hf���K]0D��<�OI�*zO9S�yʝ8�ӁJ8�9Q�ÕL9Q���p"M���7'�����F�N�5zu��ho��:߭�ti�Ѥc#F����L�[�2An��5���kq|֦<��Ly�Z���1�}n"J��D���Wì_�5|:����Wì_�5|:����Wì_��_��_��_��_��_��_��_��^�z�n�x:���u����w����W��ޯ[��[���[���[���[���[���[���[���[��_N����o%}:�J�u��������������5���5���5���5��Żqtv�������[�[� �n.�jjv�jjv�jk�jk�jk�jkzc$�錒o֦�o֦�W�Mb߭�H���|���|��f�^�3�r�����M��q5?�������rc����YG�rU�KJ��������[��exjM��%�H+���,W�xX�W�~b�~m)i����Pu��.��]:�,x9��-��K,a���`��{�w��W���m�����������&�,K�^{����0ҋb����}7�|�ȱ�z4<����R�~|� :��^�[��Al�^/�:��W���[�#I���H\5���6"ѡ�"!t):a�����k�:�.����;S;�#�􎦽�7�`M T����d���'I�R:O:��y���"�o��y���p7A`Ct7C�������/'�r�y�.��r�y�.����y�o'���y�o!� !��7x������@Cw�n��r$���"�Ct�`o0�H@Jj�BЁ�Z5B�h@�-��P� j���m�|�ρ���6�>�g��l�m�m��m�|�ρ���6�>�g��l�m�k�����<�|/_������<�|/_�b�I�Z	5�A&�h$�-�Š�X�k�K�����<�|/_������<�|/_�b�I�Z	5�A&�h$�-�Š�X�k�K�����<�|/_������<�|/_������<�|/_������<�|/_�����<�|;������<�|;��5i�Z@�V�8դ5i�Z@�V�8դr0��F5���@�#�a\� k��0q�8�\� k��+�m�x�����6�<�s�>x#G�h���<��4|�F�����5�I�n壼^�$#���(��ѭa��|���$�)��$ȟę����Ѣ��4^�F����{�/�E�h1�:x��Aćχ�J�w�ĥ���I5�H���7C\J_��Q���ҭ�1�ɮ��#���w�$����m��`ЌmMf"��y�~�Jm.5��R�ٌ�:ah��7�x�ׇ����RL;�J�K�P��6��ll�m����@ ?�ď�g�>c���7�6n�ˡ�IV%LX�1HP����S�)
X�V%��F��A��Oz�Œ�9�8?H�A�ֱ�$M�Ӷ���c	����6����0t���]Qڢ����<Ó�(�@J?�څ�cP�Lj�����>����+[-b���+[+�v����F'�щ�bzm��F'�щ�bzm��F'�щ�bzm��F'�щ�bzm��V��U���jz�Z��V��U���u�:�X�l5���X�l6φ�l�n�Dơh��-�����>o2Ѳ�-.�)�����)���)��r�X����>B'��D�]�:`�k���`�k�yʞ��T��r�N(t�R�N(t�R��GTq7����p"M���7 �#C���GQ#�:���H�[@ڽmj����@ߦ1~���c&�<4���n"Bݸ�>kSW��$���I_[���`j�u�����;�^w���Ux1ު�c�U��z����W��;�^�z�n�x:���u����w����W��ޯ[�^�z�n�x:���u����w����W��ޯ[�_u����|1���c����_�ᎿW�Я�;�_N����o%}n.�}n.�}n.�}n.�}n.�}n.��n+��n+�}:�J�u���qt>i��|ӭ$��ZH[� �n.�jjv�jjv�jk�jk�jk�jkzc$��������������������qo��֚F3z�Z��9jmk�n&�帚���wGY�91��Ɏwt��e��6�	�I_��4?�h|h���_���(�%x|�E}��&�W��[E��m
��k�rĦ�C��A�����C�̯I�<�F����F|��alU�&-�b������|�x[�?�w���Ӈ������|���g̮�\o�����|����/@��;�/�Ų,u�a�I�81X����i(�%z4��|�W������]��"��&�9-��W�u�]3q1:v�wt͡�zGS^.�����ם�o�U����d�<�GI�S�O:���RM�"�o�;�������,n����o㗓������]0���]0����O1���O1� ����������@Cw�n�� Z�ħ��Jz�C�{�Jz��mC�I�V�5�&��$�>����P�jMC�I�|	6����Z<�+G�eh�l�m��Ͳ�y�V�6����Z<�+G�eh�l�m��Ͳ�y�V�/_������<�|/_������<�|5�A&�h$�-�Š�X�k�Mb�I�Z	/_������<�|/_������<�|5�A&�h$�-�Š�X�k�Mb�I�Z	/_������<�|/_������<�|&դ	�imZ@�V�&դ	�imZ@�V�;������<�|;������<�|8դ5i�Z@�V�8դ5i�Z@�V�;��N�h��Z$�V�;��N�h��Z$�V�8�ǜ`��r0��F4����6Ҽ�W��J�$iQ��*0��F4��F�HҼ�W��Q�6x�c�r�I69y=
 �f��+
���jl��RMI`������#j�ĐB�$�I/AĐB�$�I�@��m�x	^#�	#�m)֤�6��h�Z�
-N0��6R/Tu�l
�k�i!b�b�
����yG47GZ��O_�[l�j������`y���_����@"Yz �UaH��:��y(�|�A�M�M�����H�������d���dy�nď�G�A�M[�2�_�k5ɢC��{���"�Jr�N5I"&�"4ᴀ����Rz��%&J�Z�D��i�爛�n.���]�=&�@�a�u�R4�n�A)����1)� Z����P�?j�1�|7[g�u�V�Z�ka�V����u�1=6�OM��h�Í�q�4caƌl8э�1��F'�щ�`:sX���5����ur�AܭP^��/A����u�:�X�l5���l�i�φ�P�l�F���Ly���� |4�e�e�Z6^e�e�%7]"Su�%7K�`C?,-Qt�n.�������:`�����`�k�yʞ��T��r�N(t�R�N(Tq0�GTq7����p"M��^�Da��F���G�u?����D������6ߦ1~���c7�@4����jc�I��v�$-ۈ��n"Bݸ�v�$-ۈ��`o�u����W�ꯦ;�_N�z���U}:���u����w����Wӭޯ�[�^��^��^��^�z�n�}:���u����w�)��W�~��:�_u����|1���c����_�Ꮏ|��~��;��G���������c���t+��W�Я�[�_��n|n)%|n)%|:�I�������[�[�o'�:�H�p>i֒W�N-ۋ�[�~�~�~�5;~�5;~�5;~�5;~�5;~�5;~�5:�n*v�n*F�n*Ezu���֚MM4�Z��9jgG��M���ڿ�������:��H�;�q�����~�Ѥ��O���O�8��p+���ܫ�iR���W��A^���/0x7�!ZhPrߛ�
ߑ�mM5M����|�Xϙ]:�e^��L�!p��n�_�+��X�b�Kp��%�|����*�o���2ǆ����Ӌ��:`���u_���ϙ������2�"��J�,H��-���U�ӄO��-E�iX7��ܷ�|WA�=�=0��?��0�NzF8���WL�LN����1�jt͡�,��]Q���
�o�;|���&�Y7�*��yԎ�Χt�u;���E$��wy��E��]����M�r�y�o'�r�y�.��r�y�.����y�o'���y�o! �~ ��7x������@Cw�n���$ Z�ħ��Jz��mC�I�V�5��C�I�|	5�&��$�>����P�jK�����<�|/_������<�|/_������<�+G�����Z<�+G�eh�l�^�������yz�^�������yz�k�Mb�I�Z	5�A&�h$�-�Š�X�w>�ρ�s�y��w>�ρ�s�y��k�Mb�I�Z	5�A&�h$�-�Š�X�^�D������y��w>�ρ�s�y��M��&�Ǔ`�ɰq��8�y�<�V�;������<�|;������<�|8��7�#�Z@�V�8�ǜ`��(8�J<�>�ρ�r�I��w+D��h\�#��c�(�#��F�H�x�ф��q��Z�k�����c�a P�(�
#����h��6>|/�@�LxFɀ���%�������@|�z�G+����Fb� ��$,x	G�؅6����k�����A]1|jG+���)4�9'>�2�`hi��ǓJ:5�Q�BmB�3��N޵f����rn]���ܵ9�<�9(#��� L7F
�u� �I��H�%��S�9A���ꄉ�P��GT#����b5�F��֝ӣZtkN�iǛ���y2<�L��@�#ɐ6��oy��Z�$TбJ�"<��5�4�")� M� � 85�4;��S�М.(���hpۨ+����6���Ӥ�`(غ�:C�6��`�+M�g����T��%M`;u�x6���Ji����狳\�sM�����(�Pw>�`���j��ָ���Sj��P�Pt���h��։����M�[.5kuƭn��۩�ke6�l�խ�ڵ��+[-�� |4���̴l�Ħ�Z6]"Su�%7D��(���<Ó�H��t�mWH��y�'�0�������`-,%���T.��E�D�]���R�L��=&�P�Ρ7N�����9:�Ó���6����_��H�[@ڽmj���Ө�9m��F0�jbJ���+֦$�Z��~�6�n m��@Ƒ��G[�ioQnc�Ź���;�[���nc�Ź��|��~����_G璾��'�1��?��4�t>i��|����;��LwC�����?��S�(��,Q�$���H�G�B�.�}1ު�?/��qt+�p�W�������[�o&�jn��mI�W��bߦ2�[����J��Ԋ�?$�4�t+鎒W�$��:�_Lu:���u}:Ԋ�u���RsN4�����CHI!�$4�����B�Iq�$-�� ���p+���W�������[��!�u����X��ֱoӭb߭�H�����7��7��7��54�r�[�婝�qk��qk��q6�v�mzF9��旤?���jߢ�0i+��|�qn���H>4qpد�I�W�ҥ,W�j4�4���
��/�^�,a
ѿ6�����Go��6��f����1�3:F;�.�8o��́�~���>ẘ�>|ȯC�̊�>|���9c���dC�Ǟ��o�.�/�F;�M�hoƛQ���b���<�
��0W8uD��F�_JE�Z��[���n8��~zA�	�����)��Ĭ.�f����%��wo�,�k:���Go] *i�y���Y7�*��yԎ�Τy�)'�"�y�)'�"�y�)'�"�y�w�� ��@t<�7��Cy:AC�Cy<�7��Cy+� �~ �ڂS�@9_�+� �~���A)�������-�A)����A)�������-�����> ���X�k mc��|���6���> ���&�Z$�+D��h��Z$�V�;�����Z@�V�&դ5imZH�V�&դ��i��<�V�/U�K�h��Z$�V�/U�K�h��Z$�V�/U�K�h��Z$�V�/U�N�h�J� iU�*���V�4���Z@ҫHUi�Z$�V�;��N�h��Z$�V�;��N�h��ܭw+D��h�J�iV��r�I�V�8тN4c�6�z�Q��p;�ƭ_��W�܌ M��8�ǜ`��r�I�|5ρ��(�z9 ^�	����(@Cp5���c�(�w�%��Id���"���iAė����h�#B|I�^c�� �FX��b0m�]�AyӘ���u,EūU�����:ɮy�!BS�B$�7����K�jٔ�)�l&�kף�9_�D�IX�?�-֠
�
?ʛ�~�7�Pr�i@�@���I�7�d���'�P��J²{zoS���iB�Ȝ�e����I���V��o��S�8u��@h寶��ꅵw��W�5�h��&-�6 O�H��	I, n�p7ra��7ڀ
5��ka�����#[F��l1�b5��ka�����#[F��l1�`�u��i����v<ݏ7c�ؑ�����#tN�I"��9B�!��u��F�mI6�h��b aX��Q�M	/�e:#C�R$���M�鸏��'Ќ@�:J8���m�h��(��%���Q��i]m7r1��Z4�o����t����(����k����s��s��G�e��j�������V�Z�ka�|(:KEIh� Z6j�ˌ��~�V�S`���;u6�M�[-���>��M�Z6[�Ѧ�֍2���t�-�Ih~ %�Ó�r|�ڮ���ڮ���M�!ɻ�97o�3��P.�D�Ј����9P�-t�9S�n��t�P�ru�'Q�m�����:�Ldj�mj����@ߦ1�1��ь<�Z���jbJ���7�qo��߭�ioQ�u�F���G[�[���nc�Ź��|��~ߦ;�i��?�Ɛ�����[��!n?�4~Iq��-�� ���pq�$-�����B�I8��q�H4���i�劼�xT��8���8p+���W����Ҝ�U��^�:���CH�p0~ދq�$�[���G�:�=5���*q�c����W��N����_����|1�J�c���o���Yq�bߣ�ſG�;~��qn?)Ÿ����[��qn?��������[��}�
�?��pq�$ߧZI�N��~�k�:�/鸩�qR?���?���?���+ӭ4��9n-��n-{�n-{�n-xru��H�;�a����rU��'%~Ro��D4�8\iƁn8�4hS+�p#�����B�i�
��j�x�0QZߛ\J,K�
ߑ�:���i�����1��o���%���˦�t���.�8e��`� �8��X�����#��_�m�C~Gp�-)(�!G���ǃ~o��[ �����$�FZ��Rq+�Х|���4��C�W�פ�0�M,r��u�EӬ���wH�;���ںGQ���GG�GM<�:h@o��d���'I�R:O:����`�I���`�I���`�I�y�3��] ���!������b��!��b�@9_�+� �~�����@9_�+����j	N����m��V�h�j	N����j	N��h�m��V�h�k mc��|���6���> ���X�k i��\�i_M+�I�|	5��&�Z$�>����Z@�V�8դ5i��H�|&դ��ily6<�M��&�Ǔ`�ɰq��8��Z$�V�/U�K�h��Z$�V�/U�N�h�J� >UiJ� iU�*���V�4��r�Iܭw+D���%�Iܭ^������h�'0I�<ҫHς���|� iAǜh�'1�x;�o{���iQ�V�Z�+D����8�y�<�+D��h�\�q����rБ�yޫ�P��6�/��[�6CX���!��M�AH�<��h�iII!q Dx)���ԕ����Чkw�m�6�x=0h`��u�:�B���Dִ-���n�M\f1�BY�1aԴ�8�1簺�8ZI��;�Hl:9��'e�q�\�M�T��q����j�ZԜ.���Z�&��VMPIl(CY	GE�$�0���Zh�D@����|S��H�U��Ҡ�)�ц�h]H�֏}K?sAؽ9�Z�2T�.��?rT��b�$y��A�zV�&7]��Q��	���.v~AӣZtkN�iѭ:5�F��֝ӣZtkN�iѭ:5�F��֜m���u���dm26�nǛ��y2�w�1~�A�n��`���H����Mȉ�����^;6�LCҘ��=5	��y�Y���
O��E�4/���DHB-	�� cĩ��@�o1�<���L|�n��+�Q�X�P-1)���mC�Az��F'�A�i�ke6�l��ۮ5kuƭn�խ����V�]τ��1z�L^�Sejcl�n�φ�l�n��יh�y����h�,	M����,	M�Hr�o��r|�O�"U�����!�7���97o�3�9*,e�DM�<�N��"zJ8���=&�P��q7N�����9:���hM�u^���z���ho���Lb��ǆ��$4�a&�n m��@������qG[�ioQ�u�E����;�[���nc��4_�h��W��䯣��_G琷�B�~yq�������G䒾�*u}T��8���qS���W��b����_G���+}V*�8�K~Y0��,a�4X��ȱG!b��%�,U��ZY:�o�?M0~�u~�W���W��|��H4�u8��*�-7Ŋ-7Ϛ?)Ÿ��W��b���^劼�x�*�?)�~R+���+���q�b-�����"�X�q�b-�������/�?�_4~S�h��|��N����G�;��w��#H�R#H4�u �1Ԋ��Y+ӭd�N�ҽ:�A�qoC��އ-ŽGY��7��7�^�mhru��Ɏwt��e��`�8����ߢ�1^��~��&�|����lW֤ܖ*��,g�"X�֑^j'�/�4�W��ı� ����Al��/�8�rĻ���j;~5�pq�mMg����qp@�_�7�����ٴ4�M�j;��pE�BP�����<_0u�h1�����iê"�7��ԜJ�.6�.Ɠ�+���$�AwL8����j�β��u�K�bt�c��c��hm]#���7��Q�B +| ���
�o�U���'�H�V/0Eb�RO0E$�RO0E$�<���p.� E���MA��]1���O1� �����r�j	N� �~ ����PJw��{PJw��G�l�z��{PJw��{l�z��G�X�k mc��|���6���> ���X�k i��J<҃�4���(8�J<҃�8�ǜ`��5i�Z@�V�8դ5i�Z@�V�&դ0q�8�y�<�q��8�ǜ`��0q�8�y�<�q��8�ǜ`��p8��m�F5���@�#�a\� M��h�$�0I6�k�I�`�X�z��V�$�F	&�ǜj����|4��G��ܭM���`�m$�x5�� �0�(�$k��4`��$�F	5��&�Z$ҭ��P�\�iU�Da ��H�m�O&�h�
<U��l���[�|�M�[�
�NI��NM�L&�k�J����3��t����h�Q�E��;qS5B���hO7)�`�SY�jUn)��\��;!��2��y�I9� j.ڍ�*s��G�;n�ϛAٲh �-���ro�grF�"eJ�2>jd���5���r&�<d��c^@�>�9�DiVG򰑓a��dFe0@5�	�b���H��W1���u�r�雱{L��Kb�b��5I��9 \����#ZtkN�iѭ:5�F��֝ӣZtkN�iѭ:5�F��֝Ӎ�Pn�6�L��F�#���v6ٍ�bM�e�w�1�}_�n�;�.�
���*�
���N�Z��Z��GgA;ZG+JN�16,�S�'QM*�jq�YT�mPQ5��M*� .(���ѱ�^�F�0�PJj�6�Z���b��~逧ΐ���6���^�Sj��Z���(�q�0�ܭ>^�S����1�V�6φ�l�Lm�֡h��-��(��Z��Q��7��c�Cj�D6��Cj����!�7��`-,%��D����2�t"&�r'�#z@R7N���v�D�ہru�'Q�m���F��S$o֦H4����jc�I��&�<-ۈ��j`bݩ��kqz�#��-�wx�1����w�h��|��~����_G璾��%}�J�?<��qt+���W����Á^���}
�8�餕�8X��p�W���W���W��b����_�"�
E|��)�8R+��qŽ�Ž�Ž�Žp�p�d4���iޚ��E��i��|4��4X��zX��zX���X���X��^���i_G�b�M{��h���z�
E|����N,��8Y8p�p�d4��|4��|4�z4�z����_G��+%}VJ�8���qY+��W��d���_G�"����������������1ԃH�R#H4�u"�:�J��Y+ӭ4�N��r�[�帷���:?������^�N��^�mhrc��Ɏwt��e��gN8�ÑĚ�^�9�E'�-��~o��Oo�����B�_�nX�2�^ �||���V7�оW��^����0>|7�>�`|9�JC�\,K��oțQ��&ۃ�ɶ�ߑ6��&ہb]�RĻ���8�v��R��V��x81�X�ęb���	���:�W�#x��I�-��(��cH>S+�~OJ��`?����β�`�LE�q1:F1��m�H�6����t��z�(� �ju����d�<�GI�R<���X����I<���I<�;��y� ��@t57�PCy:AC�Cy<�7��Cy+� �~ �ڂS�@9_�+� �~���A)�������-�A)��-�����-�c��|���6���V�/U�K�h��Z$�V�/U�K�h��Z$�iAǚPq�y�iAǜ`��0q�m�k����q��m�w������a\� k��r0��F5���@�#�a\� k��r0��F5���@�#W��J�$i^m+�m��q��o��m��w<�����yz�^���5��z�^����p8�\6�+Q�r����U�I�q��0I��q��Ta �F!x#G���1��F	8�ǚ�h�\�i_C�JJz��W���>��԰n�Gp4���
�m��ьOm ֘�rt	�RAka"�%���ˡp�~t;��j���p��L?|��ħ5P�I����KM�K#f[��v�X�b9Rڣ��u@e~T��mM|im��0��P5~��#S� �r@�aS�Nٺ�eJฑf�:�8�*�����T��2n�l�N��#�-յNc+a���' � �A���1V�$���� H4� �*�*�����G����c���v:ݎ�c���v:ݑ�dm�fFّ�dm�fFٍ�Pn�6�L��F�#���v6ٍ�d�v�L�O�G���y�jަ���~o_�W�ZH����lMVBu�Ubaw�RF��E��
�CZa6�[��US8+��i1�����U�_��P��u#^`)SlJ?^��څka��]0��%7D���h|�|5Z�ihP�^�*�j�v�Z�k�V�Z�k�V��~�+Z�c���Z6�C��h|���A)� ��&�ɸ�rn��b��C0t�%��D��!�7��������`�9�t�:5�7G���I�#]9�H�΢@����^�1�z�Ǜ���7�qo��4����:ޣH�z�s��-η��:�O�?���~y+���W��䯃��_B�.�x
�8�8p+�p�,W��,W��qiN4�Ҝiť:�=5"�=5"�=5!b�K"������W顧W顧W顧W顧�ѧ�ѧ�ѧ�ѧ�ѧ��mzmx��h��h��6�[^�^-��z4��z4��4X�M4X��|X�M44��zX��z4���,`��X���W������Z4�L����w,`�گ���_G�c�yb�M�b�M�b�M�b�M�b�M�b�M�c=4�c=4�Ӈ��ӎ-�-�-�-�-�-꾎)�}SJ�?7��?7��?7��?7��?7��~o[�Y7���o��o��o��o��o��o��GY��gG��Z���Z���kC��Lv������;�q����sHr?����j�$�N���LJ��C�~��n�4\5��гW�ҥ�`����iՊ�_+�U�-���������0���qm
+_�E�Ґ��k�"�k�/�5�l��6��Ö��Ö��Ñm��X�,P��^	2�z��u+�Y�W�j-ړ�[��~�������?;/L�ޘ�]����%���7I`�LE�q1<͠��6�S�u^f�ֺM��[� �ju����d�<�GI�R<���X����I<���I<���I.� E���MA� !��ˡ���ˡ�%<�bSɶ%<�Ţ��%<�bSɶ%<�Ţ��Z/�Ţ�z�w�_����Z=W�G�m��|�� n�h��Z$�V�;��N�h��Z$�V�;��N�h��Z$�q��8�ǜ`��0q�8�y�<�#�a\� k��r0��F5���@ҼHW�J� i^$+ā�x�4���@>����c�����6>����c�����HҼ�W��J�i^m+�m�x����@>����ms�m���α��<�:ǚ�X��$�x�8�n4a#J�$iQ��*0��F8�ǜ`��s�y�x5�� �0�(:#�Tc�ƌq��;��Mr�H(���C��F�_�[�^�7�(�M��;pt7��նQ�-p�H�)���h&�	59�ЁXv"hx�������M��p6=4��b�;7��3����X ����i���A�F�#s��H���s�U�zs���D�hz&�.�qB.�q����\�K&�U��f~쉰*�"v� ���
���'%l�4 i�a��	������H��~�19�� �lT���<&óBxOe�J�� ��I��vvs~��`$t�0x�v:ݎ�c���v:ݎ�c��fFّ�dm�fFّ�dm��u��i����dm2<ݏ7d�v<�L��@�/S���m2@ ?�Ǐ�Ձ�0�X��)�)�)�)�S� �(ANP�čr�u!
q:H��-������4ESQl�[;��EPh�"�h��6�M6�:MM��G]��V���[A���q �ݬ%&�r��|�*iQ������hn�>�Cu���z�0^����hZ�Z��Bְ�T����QSl9(j%A��!�:A�H"Z��r��o�6�,r"��"@���GF�e���#�:��9�6�� ����^�1�z�Ǜ���#��4����1����w�s���;��LwC��}�
�?��~I+�p�W����À�^�H�^�H�^�H�^�Hiť8ӋJq��匯�%���"���?R8~�u~�:�o��_�Ō��?oK?oE����?oK?oK_�_�_�_�_�Zk_0�ͯ�zf��=3k�����ZX��ZX���X���X���4��z4��zX��z4���,`�����w���-��������G�j�=6Ա^�Z���|���h�E��i���i������������������������
��X�M4X�M4X��б���b�B���8:+��tW��诃��_���k�-k�-k�-h��CH~o����C�hi顤?����tC���gG�u��qk���և&;Z���k�͡ɎjLs���.��4�#�Yӎ%7N8�ސ�MzC�-^�Ap�Z��h$ߡ���_9�[��拆�n46���o�� ���b�Ō#I�8U�X�W�c_���<K<�o�X�o�B�o�B�o�B�o�B��
б�����X�,`���B���$��&�W��i(���$F�аW���^���r�:�;=!h���JE��Nt��k��M/3S17��Yo�L��6�P��m]#�� Q���GM ��P󬚇�d�VM�
�t�u#��`����^`�I���`�I���`�I���@�"�jo&����@���]@����M�)���Mb�~��M�)���Mb�~�-�b�~�|;ׯ�z�h�^����m��|���N�h��Z$�V�;��N�h��Z$�V�;��N�h��Z$�#�a\� k��r0��F5���@�#�a\� k��r0��F5���@>����c�����6>����c�����6u�d�GY Q�Hu�d�GY Q�H>x�^$�� ��H>x�^$���؅�6u�d�GY Q�Hu�dGY Q�@>u�5α��6�<I�A��>x��$�G��Q�@>F���(8���@Ҿ	U��Q<҃�8�ǜj�s�y�V�� o���x:e3T�5��O�����Вw���k���%�Mi#-(�On*'Cz[I6cQ��Ҹ�۬��d�����������mD��� ΂!C��[���i���kd�M+`���8�r3"L�*�����@��x�R6�;Ȩ1��m>Z�r�����	�%l
����S��?\߫`-��MV�U�`���0P2n���^�)��.o�aPoe�oհ9�\߮o�7밫�<��{٘$t�0x���u�n�[���u�n�[�6̍�#l��26̍�#l��4kukuje�L��F�#i�#���H�$?��ڰ6�y2$��$�	&0�y���/ڨ	7bM��f@Ӎ�$8e�|ǩ� 3u�f��� l�۵��
su�q��R�!�N�o�����*��Kf��"ONm+����|JiV��(�@"y�q1 D���	E�B��z�7^��šj�hZ�>
�B��Сz�(^�
�B��Сܴ(k	Bi�P��rD��/IDk����& �%3�&�<�o0D��y��'����G[�t��� Q�uG t��y�BOI�?�y������7�qG[�ioQnu�����|����;��LwB���%}1�J�c���S����W��b����_���=5"�=5"�=5!b�K"��E�-,��_��N���W��c���E���?M0~ލ8~ޖ3�:3�:0~׋k�kE������m|�h��v�[_;j-�����ڋk�mE�����W�����������j���־a��������m|�ic���ͣN���>,�dh��4��	�08�84��pYu~b,U~wW�h�4,W�ז+�k�?k�?k�?k�?k�?kŴ?kŴZoE�ZoE�ZoE�ZoF���N���������x�x�}��U�86��pmW�ŵ���[�����n?7��~oE��׋q��o���o���GY��g@��kC��N�����c������wN?�]8�Yt��e��g�?�8�5t����E'���A����~OW���ߡ�\i�f�o�hR�����E�慚Ex	����u+�M\�5qb��x���,`��[_ǈ���m#N�<K*�,P��^����U� �W���_%�|��zԖ�hR��qf���r�:�+�g�Ot�L���`?����Ky����jf'�����S,���Yy�A�@u6�3pkD
;^�(� �ju�lR<�;|�<���"�VM@Eb�V-@Eb�V-CΒjt�P󤚇�$�\�E���a� !��ˡ���ˡ�%<�bSɶ%<�Ţ��%<�bSɶ%<�Ţ��Z/�Ţ�z�w�_����|�� i���Z$�V�;��N0q�8�y�<�q��8�ǜ`��0q�r0�܌ w#���@�#��\�i^$+ā�x�4���@ҼH� ���B��F�/��lB��F�/��lX�F�h�c�,u�E��h�֍:Ѣ�Z4^�F������:/x�����4X�F�c����y֍:ѡ�Z4<�F��h��lB�z��/Q��x|�?���A�lB�?����c�HB$|	4��7qI�Cz��Pq'��6� w>�W��yZ��T��H<�MS,O>M1�fnI��J;�z9_���h�`ַm���pZՁr��lI�nZ���ړ�I�Ǩ�M:���A���Z�j�T��.H��5E���̛��l��|�{�S��j������eʛ����\��^�#s�ᩏpC.@���cE�	d��V��B�d�݋� ��*bz&�ݦql=�7eϥ��h�O�=��3~9~9 ^�)�@=���`$x��`���GA� ���c���v:ݎ�c���v:ݑ�dm�fFّ�dm�fF٣[�#[�#S(���dm26�L��0��g�>`� ϘՁ�oS��1�T�;��w���?A~|�~|�y�w���0hI�p4<����FS�OSs�����Ss��s�t�r�+��&�$�UzP�ב�:.M��(�F�iT�[+��!�-I�$F=Bo�7�����4h��&�J�!ɻ�9>m���bеz�(^�
�B�rСܴ(w>�ρ4�Љ6�"M����5�(��9#k#�`�u�!��%3�&�<�o0D��y��'���y���t��� Q�uG t��y�BOH�zGP�rc=C��$߭M�����i7�~�o'�1�H�t>i����I_Lt���J�?��4~S����W��b�Md��ґ^��_�!b�M�+��ӫ��b���ӫ��b���c��Ӿt�c��c�趾s�c>s�c>s�c>s�c>s���v�[_;Z��������������������������������������������-���[_;j������ڋk�kE�����ѧ��l���mR��E���>,�a���(����Bb+H��t�X��8�_9-�1p�ߘ�K|��5oʹ�������Q�|�Ӈ�hӾv�i��i�;j-���qi�qi��i�qi�w�ז(�ז(�ז(�ז+�kU�鵪���U|zm��=6�_�j��M�|צڋq����z-���[�����n?5��?5��?5���:+��Lv�91���c��юjF9�91�AɎwzF9�ӏ�N?�]0�izC�Y��7�?�×�LB�H9���Z	?����_9��_9��_9�9��N8,ƐаJ2E_Te��M��M��
�u+�uX4�B�i����KF�,a�^	5|z���/��^+�ЮW���_%�-U�iq"�n��0�>n]8|lt����C�zd�u�����X��H�&��M�jf!�Yo�L��ڙd@u6���y��Z Q���GM ��P�`���y���o���"�j+�"�j+�"�jt�P󤚇�$�<�&�"�m�.���kn���]@���]�)���M�)��-�)���M�)��-�b�~�-��ýz�w�� i��m��|���N�h��y�<�q��8�ǜ`��0q�8�y�<�F;���a�@�#�a\�k��+ā�x�4� ����x�G��Q�@!x��^#b�؅�6!x��^#b�؅�6,u�E��h�֍:Ѣ�Z4X�F�h�c�t^�<E��c�tX�<E�h��?�C��Ы�u�B��hU֍
�ѡWX؅���ޣ�����6>����c��؅�6u�����HX�>�q��y��`� iAǜj�����
+@ � �:�f�S�@����HyXִAޭ���鶦KH6�i$�rַ^��94�#`dڍ~R%6�
Z����sA��i�&�#�*c�1�~䩺�m�	P��5�0MmS�D�0��t����Ff�m	��b���6�r6����de��7[h{3{G\��x�E�U�e����U�e����"��CU9�¯c-��������� �ڮiSߘ������ ��.��r �=��g��^�_E1�S ��� ���7\@�D@�D6|�!���jd��������fFَ�d�� j�?\H���n��26�٣[4kfHݍ�H�V��tK����F
��TO#�闫v$Ӊ4���;��Lc�1�T�=S�Lc���?�O�����t �-D�*\�*\�j�F�A��[pRE9HEYVBtМ�E;�ea�Hzz�JL��Z/چЧo����נ�����;�ګաCPC#y�th�":������9��u5��v���o�8غu5��ֹn�I�HX7At�t͠�]:����6�<�� Du�yѮ��6X(���pt�P�:����$.�%zu���oӭЯN�@�1��c����o����|���|X�M4X��zX���4���X��Z4���M4��z4��诊�4���|-Å!b�M�Ӈ�{��A��Cjߘ�ږ0�־`>6�0�ַ�86��.6���������l�#K�ͤ�-��i|��Y,`��ߍ�&��.E�>,�*�mU�鵥�m#W���"�|�v�ƃ�[Ie�#i1?���4�����Q�/�Q�����2�O�jF���A0�����u5C�����/����h�N��ir��,�Ġ1n-�\1%�%�4&%�%�h�bW���|�i�|�|m|�|mo��0��󶥊�U�_�����x�����R�|�ux|�|�U}W��}W��|�Ux���������n���8��Hqk[�k[�kU��ګ���W��j���k�1�A��ںs��t�[j����5=#��s��1�!��VGk�	o�Z)/L����JOHq/L�U�]^��f�j�\Y�!qfߣCn��IJ-�J�[����jN%|7���7��o5�o��Q+��W��D��gR�U��u>k�J3H߭Ij�Z���
P�\mÐ��C��9͏HZ4��I��$'H~)<��1�:ɯ3q���j je7����1e�1�wj���nי�5��t��z�7��Q�O2��y�v��y���o���"�jjF�"�j+�"�j+�"�m�jv�"�m�.���kn��r�j.�ؔ�m�O&�h�k���h�k��ؔ�m�O&�h�k���h�^���ýz�w�_���޽|;�jתmZ�w�������n�p7p8�ƌq��h�&��<�<��#\�$<I�A��l|�?�����H*�8F 0�L�F�#�Ě�j�*�#m�t����������B� 	��Cδhy֍:ѯ�u�p���ЪL��I��#�W	hA|��©2�����$aWX���F�"+n �LL:�-8GC������x�χx�|P,_8�ǟęXS�Σ�l|tc��h��Gt]bb�� �Z<�>�g��^�V�G5:Ʃ�W+ɳM	�)�L�-��Ĥ�|�! AZ�jO���H��j֎#���&��b�F�4��rrH�D�*I�0v�6$M���*{���Lvbc��l?[��ku��{�>����r�9� ���M���7sDF�2:�JT��誂=�	  ��R'1Lr���>�c�=9��l=�`����������[G��ӆ]����������������c.@=����`�sױ�t���{G\�e�TDTCg�� H~�je�n�ϐ$?`�vFّ�c��!�ϐ?\<�hz�w�%w�%0T@~�kf6�L��H�g�z�Pz�ަ�����A��A��A��A��A��A����Ǫc��L`�c��z�ާ����}y�kEH8
�_�����m�Qt\w �$EIV%LX�T�t��F�#l&�BK��j�.:��o;����"��z����7���6�4j��&�|6Ģ7H
HX7��8��a�PC#w+K[a��joUz�W�p$k	EI��SXJ*M���a�XC#GZ���5��jk�婯�;qy+ӭЯG���+n)��p?��4�����B�~S�!�H����[�!�W�E}�O�?7���R#H4���_��_����di��Ա��R��hӾvԱGh��q�Q�|��hӾvԱGh��qmjGw��IX[ CK�A2`�A2c�A2c~0�9��MʌS�R4�h�bt�wx�
�p����@DߌK,a����R&�eF�4&$,S|�i,�(�mW���W���4�H�Xͤ�X�A�ӏ�'��<��+�*��a����x8+��]m�����r�nZj���:�Oo9-(�?$���7��u���-6��.�0'$,Bʌ5o�h13�;�*�mU�?mK>;�h�iʌ5d Ѡ�ߣ�z�G�Ҿ������H8:+��mW�hگ������Z-Ãh�ZѤ?[�kU��ګ���W��j�G�����c��9�ںs��C��91�OH�;�#���sHr?���Ě�$�N�8pNt�I�'N×�^�=�F��)��|ܷ��ko���4�Ř�w�jJQ�Ԕ���R/��R/��R/��R"���3H��D���Hp"@[��#~�%��jK �\m�8�tねӾu3����_�ސ�h^�]��$'�&<��1�n#W���DL� je7����1e�m������mj���nh�Gk�&�޼�:i�Q�O2��y�v��y�� Ed ���PCR5�PX��PX��lCS��XCt5�7CXCt5�ClJy6ħ�lJy5�E�X�_��E����m�O&�h�k���h�^���ýz�w�կU��޽|;�jתmZ�w�������n�p7p8�ƌq��h�&��<�<���\�$k�$�� ��H>����c��؅�6>x��#b�Y ��/�?���{�H^�/�Z���F�:Ѣ���A\PF��a�Z5�p������:I��RdaT�1xDW?�3c�LX�#�GE����&W���5�C�>z��`�U�:V�dn壠F�"^�AD��\P�-��2&�H�
� އ��1Z�i^w ��/ m���(Jw��@U֍q�T�1�ڻ��j./M�z�:���}:�I�n[V��xZ�;^�!V��u)#���P)5����/r6���� �-}#[D�j�0�@�M�pkM�����0��������`i�+U�|�n��ov�M��~�CZ������9�i�S�]�A#� b >�D�)�b��] C9�ӟ����*�+���5����vG�����C.��H�H�H�H�H�H�H��a�=���G�3� ^c���1tO�:~�4�d��"nț�&�|����$M�vF�?b4���CũRH�u����Aq�uíؓU&���>`���G�#����7���-A~Z�ȩ��s��s���j��j�$�A��@I��ժ���_�]��$}S�i#zHݎF�A��[y]AE�Ep	�%9mN[X�1HP�|D��F�5.p7cRK��G|����b�������,C���&քmp9S\P�V�&ե�r���D�'Lu��B����]n�I�5�B�������Q�څ��Qǝ&��g{�:�A���zG[�ӷ@���OI���3qt'[�Ә�!u�;�~�ۋ�9���8Y>h�׍;�mK>5>hp޾h�׍8~j|�R+7�Q���ä���2�A~0�1� B�����jF'��������ľD�mQ���~M#�|4����W�z�>sQb��l��V��!����k�[�t�I;�#���@uԘZ���)Yh&�ȟ5_�Ɛ�ּ�:�[�-�bB�!mm%1�����Gz�]f��O|�W`��}|�Wf��(��]���D!��J�L��B{|Qчr��+��T�kW:��/��c_,��C)�1�OÉ�����0�
��$�Ҿ����bp�@�����Z5#��_E�Qcg���������J��͢��������U�_���_���Z5>k�mE�pmo�ŵW��GS~�&���*�;��������;�&9���w�?�Ó���N?�C������r8�]1�St��49J�Z�/L�0k��Hq?������]^��f�|���|��z)��pn[�pnF���B�ͿF�ݿF��i5%(�HhX!�`-ڒ�^�	���pm��|�_9�Ӿu3�́�~lt����@�����q!:C�I������7�����L���a�Yŗ���f�jj���n��׈v��n�̣��e4�(駙�oDЀ"�VMAH�ԍAH�ԍ@Eb�V-�N���N�RMa����S�zJp/IN��ЛZ:kGC���w>I���6�t&֎�s���|<�j���Z�q�W�7����z��V�Z�+@�Pq&�I�iAĚPq&�H|�#������(� <I�A��l|��F�/��x^�
<������?��*�$|$�η��|@#I�C���L�$�ѡ5q�p�$�4�4F�F��hЂ�t �/Dk�7� �/
��0��L<��H���0�A�^>M#T:�0?�������_�]cm+��^#\j����7
/����1�T�\5��u�@|8�D�&H4+
ǀ��
�^��xx��1��
��M��0rjF���M���N��y�R�8�N���w���֑��jb���kU�&�-P�V�	��<�텯�� [/v���买�������L0֘j`D�n��=ۯ��*��<85@A��?s@�<�By��dI��a�H�� �O��>�D�)�B���@��o�'��
��������o����=��2��������{s��e���S �h�/}��C���H���&쉻l��16�M�l�O�F�#L��H�$i�4���O�t�RX��:ˏ�F�W�M�yj����&���>�H�����V<Տ5c�X����f0`� ���0��݋�ˡ2�L�)#����>A�|��ݎ�v<�/#ȶ�-�
.�����-��jr�H�9B&�MQЍSZF��;1�#�`�*|����P��k��]:��Lc���SS��S���O!t�p/IC�p9R��F鎠7L���1 ��6��u:M�I�m m��z�M�X57x��W��q_�GS԰1����N�����/�Y&:����Qb���U|J���U}�U|ͯ��ͪ�~Mu~m|�R+>aF�0�bG��l��β ��FZ�@�ȍ|Zu��ů���J,ֆ(���M�95��)n"!�XHa�"8u�<��C��hb�RQ�9+C���pl�4�К���	mkB��8�5���g㨤yhS������KD�7{����;�m�&t�W[^�i����e�ڌu�K�����r�\�5F�:�TO�R��S�Թ�mA�mAj<�1x�6���0M�\�-��F!$:,Ht.4��R�Ɨ��bs��Bic�%x|����.����?,��;��;��jA��i��Ɛpwo���ߣ�e^�ŗ�?����YC�e^�ŕz?_��wLsS�1��,�!�����`�LN��)�qĤ�E����N�8�a��X�Ǥ���I��;�'�"ѡ�+��W�p�?;!���>u3�|�gN��Ν󩃐��C����7�,��|�_;n�s[�ۗ���Ι_���h�.��C�zd�L����������O0�L䶠�&��L@��mA�Vm�A��mv���Sj :�V�Gk[e�(�x�Gk�e4�(� �[� E4 ���PCR55#PCR6Õ�l9X��5;lCS��5;lCS����X9I/G/%���%8��mh�M�	�����y;�'s���|<�χ����q�W�5j�ƭ_�������+@��h\�iAĚPq&�H|�#�����0x|�#�� ���(� �F�hQ��
:���A{��X�$:�����<@��y�q��C�ʐF�w�c�ǈ�&�/_�� Ax:W�#�WX؍&��ѡ��Ax:^��7�|F#W�����y|DHR�5q@U|:#W�M� Z,x���U PV��P��m�Z�7��F�$
�	��DP,u�5�����#C���_�$�z�xwG	��ヨ��c�[B��ؒAf�|ʞ!3B�;-\�n�$i�7r�'^Bc.�&�Iy�t�l�0{�Q�W�CbT؟�J���?ƫ��v��l582o�'D�{\� ���?{@��R`6@1��PPON~������� �;0��sU�SLB��� ��t�"}��S��r~A�R'�H�E"}�7��������=�1�R'�H�#�	�}vG�G�G�G�G�G�G�G�? �	����� �E1���S�N-��s{<	�qCNPӔ4�8�f&ى�bm�bi�� :~�t�bi�� :~�|�l�p�k@k@����"C�<��/Ȓ��/ʚ����	ǚ�"��f��j����?��GS f0`� �`f-���7c���?�/$ˡ1Bb����:��UΆ�'CU�ݎ�v<����N[IRF���$oX���*D�(\׎�6��M�5Z':Z��܊M�� �7��6��#RV(��1y)��7�6�`W����H�Y�3�zC$q��ǜ��|;�$m��@�OR��_�2����{�u=^�qS����W�~֍8�wq����G�rc�1��t����QޡEj4�0$"��l?Y��T���6^�a�о07������F6�ɥŵ�ST�ҭ5_�+MW_|����,օ�>,!��F��{���o�m�j�LQ��pD���:\'H9ޭ,���ц��yZYc��u�����,փU�9H�O~jfǰ)�����5"^5�c}i�R��M"W/Ӌƴ��Xޮ_5��&"�Bk�0�]i.�1��8M�\&Ԩ�R89�R��A\tA�ִ����Z`y��t��ܱ�H�������4��P���8��	�M>E&��18���ӇƑ��%���J���J���O�-_4Z,�w�YA�ݿG~�&%z?���bW�����LJ�~,�����槤c��8�YG�r?��#�.������鈃�h.��?����NG�8���Ą郁�zawN-]0�zJ�$鞙=�=2{��HZ4:`����W�gL��ΜZ6:qh������=3��zf�t8'���<]E��o�	��$'H~)<��8@?�ڃ���֠�+51Y�m�ٴZ��wm��SP��Cp6��;Z�(�kP:5 S�̣�� V�@o� V������i�!�ͱ�m�*F���kk���kk���^�RK��Iz9I&�N�)��%8kGBmh�M�	�����y;�'s���V��j���Z�q�W�5j��w������iQ�V��ң�*1�ң����>x�"C�Q�$x�"B����<!�^#b��4^�F����� ��H,�d����
�ޢ4���t4�����Ƅ�4F�w��� �����Aޡ��Ax:u��$�4�4F�F�����Ax:�/�ޅ�о#ca���y�@�$�ޅa Y FV#Dn ��l�F�^/ �LI_��A����ޏ�S��J�#���$
���~C'>��Րu�jn!����&7HZi&ĲQ!�ʈeq1qZړ�C�Z�ޱ7�I���r	k��
T��4���b���b<n��nn�7v@MmQ��6�	���b9����f�"j�4ݩᭀ˖�.N~T�������vDZ���Ƙ&6ض��r~�?\�\�1�5@��Lvce����� ��t�"{~c�f9b���1���L}��L}��L}��Lv~\�)�>�`$x!PB���aWaWaWaWaWaWaWaU�I��TU-�A��y<�7�s��#�nǝ���SbTؔ4�8�f&ى�dM�7XF����$i��i����Di�7X:~��1&�M�nѩ������I]�g��M��OS�f脍��Z��+ԉ(BQ�C��ڬ$>�@��0c���0��.����0�ϫ�������/��_���?A~~���S�����D�j�y5o&�~}_�]�t��ռ��V�7�k"�&��5�h�����$EU!�bշ�����'	/懔$6:+�J9Ԧl�	�h�<�@����p���:I�jm�r< :���Sw�s$�G ��O����n-&�����L�-ޙ�i�rc�e�x	���Б[���L�\����7���k�å�����F��w�MW�k%�����mjӺCJ'�e0�51j�����k����kn��&%!�����d�,F��b�Lx��Ҳ sJ̆NJJ�Q)$2Yš5(䚕ZShx�8[Z����AIi�5V7�^5��&ԯ��c�kK����i�Q��A�D�:._6�\%�*��r��h^5���zUq���2�6�<!�r�z����;���\&ԫB���[M�7p�N4��K��A�����i�![C�K��~E�-��L[Ecb�
�������U�_���_����,�w�YA��i��M-�8�U��bW��i��LJ�~,�����s��1���4�s��ڙd]:�"��5zC�1�%!t~&91��d��?���L,␺8���Ą郁��������4�A���C��za"�Z'�L�X=3@�8����.�&��~'��H�BE��o��]��O0�Ly��`��'595�1ɭ��5m���l�-�h4��Q��:�M��jk�j�7kl�����ֵ�V����)�@o� V�@o���d���؆�6�6��!��ab��-ab�����z9S�G)%��$�%8d�l��w-	���6�t&֎�s���|<�j���Z�q�W�5j��w������ң�*1�ң�*1�ң�*1�>x�� aG��Q�$x�"AG��Q�$!�_�����@/u����� �������Ac����?�� c�x&��ޯBL�t+������n��Q��'���J�y�h�c��F�F�$��	 �&��Ѣ4�4 �/B�ס\:I��5q �$p�����?q\.��48�������jmɸuZ��K�٤vCY���a��Mc�����H: ��!HP��s:�lѫq%������F��ީ��́�l���ď��[��ն6�O��M�Su��1:�{�=����-r�'I��n�b�ݺ�?Oa��1��G��(?*l�\�~A��?{�90�AQ�&�$�U��7���U�U�3�[ ��V�*��l��=�D�)���1�5l9��rrr��L}�: ��v����b��)�o�aWaPOױWaWaWaWaWaWaWaWaV˒V�a�䕰�И�e��y9�a�*{��'րA�{~aR��BPؔ6"m66P"l�F�D&�ae�����H��C����(	��:~��1&쉻n��@�D<n�x��!&�MT��@ >��^�G��Z ��*z�*7Dn���A�o_�k�z���7���#z���-��]巩��oz�ަ�y��`������ո�ջϮ�tOS�OS�N��/Ϫsz���ͣ���$EU��baY�ޑ�mF�7�Sh�6�i�[6�I�{�q-i�.��ۨ�yZK �?�ڃ��fѤ�ͯ�8Y���7 4�Dm�9F��#n� �&�?�C����r���9Q(�mo���Z�Ҝ�SD��!�U����Ĥ�j������k�m�m��W�ݏU�mc���ͬx����݊�@9��ԉ�j�[T&�ŵA�wb�������7�Y� �5��5ĢrWY��1"%�>���6�a�r�����s[^5�s[V5�{oU���oj���T�oW+օ�^�\ޥH7�ø�a�Xm2�6�VL��R��Ժ��q�b~x��A#
��%�O� r˰9Y�\ֿ/P�$a��ZVb�5#�T��p��M_E���a��0X$����ߘ~V,KR'>`h�`h�`h�h�S,P�����������Y�E��F!�F�piA�Y�GK~�&��M#H84�'�YW��e��p��;�&9��f'Nc�K�bN�K:�Ł�SLr[��Ł�L,rc�?��!�����q`8��Ą.�$"�8����M�q!7��.��໤] �� �����G�?�E��.���t���.��฀�'rsPc�Z���cV����Y��:�-�h4�͠��F%�p,����k�j�(�kl���`�k �{P:6�;z �� +|�<�&��Y6�6��!�ͱ�k+&���kk��N��ף�:�r�^�RI�S�6Jp&�Nr���Z:kGBmh�w>N�����y8ի��~�V���w{\�k���*1�ң����>x�� c���x�"AG����<!�_������</u��d�Y ��6,u�Cδhy�:u�Cδhy�6u��\$7	 A&<#�C�0����D֪zE%D�ԙ#q'�=	4h���zh�c��&����n����� �$8I��5�I�^��4,�F����ܛ��c���F�͹R0��C	6Tg��,�I�_]d�7����,�F�/;rTORt�P6�R�䣭T�'B8ԑQ�H�M'�4�thb��=�P��pQ7�M䠤.n�l��:�*O\|�ƫ���(ODT��a��{�6Q��r{�S؞
�0vTD�S�MnH����{��m7;M�~�0v\n	��)Rc�Bc����kT�:F�\Z���`���*�*�)��9bsݲ
�l������A���o�s~�������7��*�*�*����S� �1b�O�p���s�lU����}vvvvvvvvl�%j�۫g����.IS��6���{ ��TR<�BT�(lD�li����uu�M�M�S44�."l�&َ��?D�>@���x�p��#BF
���i���$n��F�٣[4je�@�1"b!������T���T�Z��y5o&��ռ���
���(�J eWym�az����k�I\���oy]��{Up��3���_�]Z�²0��)���M�B5GB5I�&��B�!R�B吚&����A�"��k#鴪w�D咩,��oN��Wή ^�3����|��Q�L 
K\J+IF����C���m��էzЬ����Y��7Y��5Rm��m���M���M��M�[k����xo����ԉ�ڠ�kn���mP,�x�<MW������moT�ǁݏ���i�
h�Q#
Ȟ&&:�T���&�i����4�:�T	�M��M-
åXנ�kQ/������	�󬲕�YJ�:"WZ�i�zЬMW5�U�A��ʉ�8�oO-N�	i��bL�)&Y~_�:��+�R;���Y�;�u������e�VN���&�7����b}FA�@>A�d׵i���SV�0|R�(�<�6�����m	��4�\&�8�5q�jX���^9M^9M�E��F'��B�84�p��-ÃH�LCHq1>k�+ �үG����!ɎwLs��:�OH�1�Y���f�I��]&�io��j�d���&:a����r[1�e��N,�p�?���Ą郁`�!����'H~)7�Ą��໤��E��,k���~���4]����G����~�Y-�:�m��5m���lu�Z��Sk�KP�M-a�bj�Pu�f�Yk�j�M���ֵ�V����`�j �F��oD;z ��Cβju�lCo�b|���r�kk��N��ף�:�r�^�T���I6Jp&�N�)��Z:�GC�h�q�N7á��y5�ד\�_��ד\�_������ң�*1�>x�� c���>x�G��Q����b����<!�_�����@/u��d�ر�6p���hЫ�t*�F�]hЫ�l*��Hn ������0��~c��f�l~XKQ0r����F��	 �L�*�zh�c��F� �H��M&<I�>N�"L������%����6�8F�j#P{�aMm��GS�HD�Tܵ��#�ݾ(���r����e���kS��E��ՑB�7���Q�u��ƪ��u��H�o�詃���?s�("O~�V�6F'#�����(O\P����L}��OӐl����i��~���͠MmQri����m��.v�)�������I��7_�n�[���I��O(*j��l�����rO~bpdߘ�
�i��V߮Oհ>�__�A�ᭀ�ݦ�P{��������c�����e<R	ª��b�o�g��=�U�U�U�U�U�U�U�U���@ce�*����-73�`PvJ��� 2���	��	j��BT�aSa�M�SbP�`�e6�M�Dg�O��.$j�"n��$?`��g���n���ϐ$?aU���#Cg�#S$m�fHݒ7d���dm26�L`��H��>c�����/ڨ/ڷ�R"�/ʫ��<�/#
�޿7�ڷ���at^F��V�?��Hq&��y5n��0��
�¤-�k"�7�&�&�7�7�7�t��l:Z�65�lkH��ԍ�Ge�و�b$�F�e:%�i�*0�d�K8%�F��c�D�F�i��;�m�|m����b��b��b��b��bM�bM��������[��xo��m`������8M�p��k���k���k50�50�;�����w�W���4��4��4�FW<M-KC���j\�mQ/��/��+���Q7����\�k�:���ƵR��T�kU+�JƵ�Dִ+����⹯2�kL��Ն����b���mF+�Q��R:�Ԏ�m_��qI3�������;�u�_]e��Ye��Y}x�\�&�7����isx�\ц�da��ZV�,��Q����5��D�`V��c[���!ӳ~@��[*04[F�c�"�
B�m!rāJ���*���cN8[�	m�����j�-E��jM�گLrȷJ���Ƣ�����b,cS���t�4�9X�1�n��So�9-�1����!91����%�#��rX�c����Ko�9-��n��Kt��[�?��!����� �Kt�rp��'��P?��!�D������"y�r��'5�Lj�51�P�ƭ��Sm��Y�jef��4�͠��7ըQ�V�GmZ��m��� ��<�kP�@�j �{l�g��m�v������i�����i����"�"�^�T���6CX��k�)��%8d��h�M����ܴw��&���
����
1�,��Wá�V���
1�!F;���xQ��
< �/!�HB��]��
�^�w��.�{��/���B���Q��
�	��~/�W�����y�@�#���A�Fp���aWX�iZ�_�A�� ���$��7�hrLY6$��qZ��	��!��Q/�'� �_��3^4-L� Mԍ����+?�D��$�!�#�3tpF,G�i��W���5)���;Y�΁I0�h��rۼ�<ݒ6d�����&ٔ4�M�bF�P��J���90���s�\�L0ra����s�\�Wd�X~
��j� |���Tǻt��l��\�l�����dF�k��>�1��{�>�~�1ٍ7�`��{A=����Pl=��������q���dM�dM��I�lN[r~�
����V�V�V�\�\��h�aW7됫��<5<5<58����s~��\�1�S�1�S���.�/���.®o� �r �������#܀.NО�y=��{��������4'h[{T	�p'���*{��>`�0O��KT%��ĩ�(i����6�M�Dg����.>\H~�C�������$?a!�	�@�D6|�!����	* j�$?`�v:ݒ7d���dm26�L�&0I1�I�?@� 3��ȗ�T�/�X�-c�����:X�-c���i�4����>�������/ϯ&��ռ�����oy�F�9��S��%Lo�o�M	�M	�o�o�o���(��ta�M�B+^Fƴ��i��GP6��䒘ܘ=+��۩+�O��,�p&%|j��ZY�7Yf�11�iD�4�/�/�/�/�:�TN�����ԉ�mc�������mo��mom���&�8[[����[����[������x9�w������,��+��x���,��,�xU?�-�Y��h^6��������A�tb@�ăZ� תH5�MkB��hQ5��i�Q��J�kҺ�ӎ����]Xm.�6�VK��Q���b�Ԏ�5#��W��2��xj�,��K/n�'Ye��Y}����'g����isx�\�&�7����isx�\ц�da�؆Ll>�h��'����	��c���pZ�^����͢�����������_�U��Ż�+(�M|�R&0�MW�h�-��_��c>q��1�/��1?����f ��;�#�^�#W��ɭ��4�����7H�)��95�1����βs�:����KN�[�1�b�Ko�9-���H%�C�-��n��Kt��[�?��!����H�'5Ę��&�!��?��c� 1��A�Kk�լjcV���[c��52�XcZ���6�KP���B�ڼ�;j�(�
mm��֡�kZǝ�j �{Xk�g��y΍��ަ�t�XM&�t�m�M&�t���/B*D�b�!�Sd5�l��M��I�S�ܴt;���r���|<�χ����+^B�w@��,F<���Q�
>O���!F;�(�x�����G���$!x�^ b��^�_��+���/u�C��!{�H<�
�H�1���HB�w��Qc�^�z����&�z�вL�Fu��A��xHF: �&��֤�G���KlM�'A�a51�M;��X�'w��$ă�Z`U�����%���JH-@�E�Et�R[���c��F�4�BKE7�����S�0��sL���	�t����>nؖ�eM�6Z�-P�'0�9�	�0Na�s��W9���|�j�ڮs�i��j�ڮ�>�1��>}a�*cݺ�L{��a��	��7A1�	���9�>s\���L��L}@��c�0�kL�	�a�a��)�lP�e�Rb�����M��J �O{bp
�k�����sG�����h�4{�=��sG�
�
��1m��o�[~c��9�c��9�c��9�c��9�c�=�dx"�їd{��9? ��=��/ ^	��ڤ�M	���4-��[{T����� ���=��{G\ b#t�t�:`�0O�'�T%��ġ���(& F~�������u�TD��F�Q��C�5Q� j�>@l�� 2ր2ց�u�g��h��52�L��F�#i����v$��$�	&0� 3� ��z�Pz�ަ�y�~Z�AkH$�$�<�+�{���>�ϯ#zH����!�9B��j'A�F��V�7���rڜ��*bĩ�B��7�&��7�7�7�v�N�	��;zQoJ-��Ekȭy�#cZFƴ�m��v�Nw"��!w��R"W�<Jc���J灥�f�,�+��V����mo��mh�Uj�W���;�&���x��U�j�MW���5]f���u���U�j��WY��;��wc��ǁݏ��9����w���	ݎ�'tN���Y���y�jJ�mO$�S��kB��T�kQ(��Mz	�rA�T�kZMkC��y�m<�kN:�ӎ��㩭8�6�VK���ͨ�sj1\ڌ_�ׇqK�Pe�2L�&w �;�I��:�/��������1;?�N�K�����19#
��²r0���)��
khڴ���)��I��Z{�j��4�# �&��P�Y�`��u��%`؁�����
�����Ӎ"ćN��Ų�F�\%���)�j�4���)���%�0�w�W�~LOL��G��Jn�q4�'�Vo�9��1�O1�iy�����+<�95�1ɮ�q%��L�.�2h��ɭ���[�S&��L� n$�ٸ�Z����d���%�Y-�:�mA�Ky��[�u��f�Nm��9�n$��R���%��Ě�7kP�ƭCS��L��52�Pc�f�im�A��m���6�cpmZ��k�j�M����Z���k �zl
ׯ@��
ޯ@���M&�t�m�M;�i�pE�w[�pE�q��N2��JR;�JG�b�-r���-+��Ҿ7á�|:�ǐ��/t� �1�F:���:�B�w��P���x=D/1�B��@�η�y��:��W��<�z�_�A���U�<�$ѯ��H<�z�c�W���x���0��l �
�G���Mu_���r�?��@u�оy=	5 u֚Q5�ebڸ��%ѡp4�p3�3A�������Ҏ�
�6�b��$ҫHׂx�����Њ@ؕ�E�Jp�j%9�$ռ�����u>D�*N�\��s�9�tݱ0l0�>`��������v����7rcU�|�?}�=��O�O�X~�>v�]�j� |���Tǻt��n��@[�'��|	U�rc�0Ll=�/�&9�Ls\�� �ݦ	��dM0LPOPi�b�j�j�jp
{���.j��M
 �P�{��V�V�\��O�4{�=��sG�����h�4{�=�S�1�Sߐ[~Am�d{�=��vG�#ݑ���їѐE�������c��;? �)�c ��G�? �s��@9 \��dN��;? �����D����[�V���t�t�>`�0O�6%M�CM�6	�XD���!��Cŭ���Fّ�d��7\Z�@�D6|����랥G��G��5Q������526�L��I���y�L`�c�~�� g�>��oS{���*A$P�N&�N&��@]�F�X��tW�Z��t\�:�M#L���)ʗ:.����0��jrڜ��-�J��*bȩ�"�7�7�7�v�N�(��)��h�މ��9�NבZ�+^EkH�i�F�kH�הN��NS����N�R;��q|jhI��<LL4�hS��l|o��Zw�N�sU��-��m�7�f�,�����o��v?���o��v?�����;��wc��ǁݏ��v<����;��wb�ZL�I��I���-�C��hI���&��6��M�<�6�+��
ƵR��T�kU(�օZ��6�uO:�����Ua�ʰ�eXm2�6�W6�ͨ��|jG_��Ƥt�e�&Y~I��8K/n�۬�	�b�1x�\�&�7����isx��g$aY9VN)�����Ʃ��T�q�p8�9�5N|S�'�r��К�C&6 �&��Ll��d�k��Ď�kO$ͩ[�I8F�y!�I�0鬱!+���b�Ɓn���H?%�h|L|���߯L�雉e_C຾��u}����_��0�St�sP���]!����H4��9�@c�DYX@u��f�5t��M�1����5�Q�5j�լjcV���Z����d���%�Y-�:�mA�Ky��[�u�׭���Ķ٩����Lj�[l�I�cS�Lb�lc�f�Vm��Y�jefٴ[f�ik�Xu���ڵ���k�j�7�z��W�9�6k�`V�6k�`V��o]�V��o\o:i��o:i�CM;�i�pE�q��N2ɮ�ĥ#���k�
v��k�
v���iU�&������ ��~!V��ǐ��iU�!{�~�5�G �����G��B��@�/1{�H^�:ޡ�[�*�z�_�AW��U�$x��#�C�l^�yQ�VҬF�K� ���I������w�`a���p�B�� ���m$�qčk�gq��(�JU9s���Mj��°5�qJ�}%Ȝc�4�H�J#��cP�����szٔѫ��$��2��-}�
)�n�"I����*v�����S��s�U9�
�*������W+U�|�>s�9Ϝ����j`+u��n��=����i���X|���Tǻt��i�Zo��kt������4�1��Pi�cu�u�L�T Z`��}A�	� )� -��p
�j�j�jp
{���n˓�؜�����r~�
�������������h�!Lr�!L[~Am�d{�=��vG�#ݑ���ѐE��������#��0=�dx����������>�c�>�`$x$x$t������Qɻ���`�0r�-�S�����R��BP؉��&�ae6�"4��Z	���"m��fF�$j�-h$j�F� �>@��PBW���"��
�ϐ>@�����L��I�F�m26�nǛ�$�	&0� 3�	D��m[�޿-A�T�$T�NP��$�t�"<�*\�0A$Z�bP�dDy�t .�$8�#hX��S�"S�"S�"I1$TŉS%LX�T�U9UNUM	�M	�M1���u�E4Uo�m蝽��s��"��V��֑�Tj#h�iyA6�בZ�9X���8I�Y�������C'%n#$2Z!�5PՋB�Zi�����w�M5i��1U�*��F��b�Ta��11bb0��a��&&?�����;��wc���	ݏ�R'	��b��b��b�D�mQ/UI6��Lڕ�ڜ_6�WͪU�j�|ڥ_6�]F�Σi�Q��8�kN+�U��*�i�sj]\ڗ_��Ƥu�|jG^�/�gp	3�Y���	�b�1�__������isx��g$aY9VN)������i��4��5��&������|[�ka�KP|��5���9�5[ZS������mhSrZ]�& Bs�䤶�+ u��DKa���E!n.��F6>a�Y�dF�|�гp��[_%3�����A��&/L��Â[����So㉉��&&�8����bt��ˤ?�^c����bf'I���&�St��L@��b�Sj�M�n%6���קX�zu�W�X�zu�[c�j�cV����X�zcצ1M�jcVٸ�DĚ�51�l��ͳS+51Y�1�ͳh4��1e�1�-ch;�����6��m�6���ڦΣjl�6���Z�nk�Gk�j;^�QΎ5��[ָ
޵�V��y�M+Κq��q4���1�|���q)d��Mq)dҭ����|�X��p��$V��*� �$!V���{J�I�+�{�~ҫRAT��Ь$k�
q{�~/x�ŏ�x���?���[�<�z��oP��H<�?ă���x*��G�o���xXJp�`mI\�	���B1���υ#iH#Dn����$b����9�ܜam�wp%�
őDP�4�DCj��c"�5��
�Ќ
Rw=53�D��nՄ����Yޥ���{b�?Aޘ�m����&�$nѭ�5�L�6X&�(N�'�-[@�m��F�Ȍ���O�O5\�W)���|�?}����g���t��l��@[�-��u�����f&;1��i��T��V����{@��q��� T [ll��l��l=�9����e�L	�������� ���9
�
��182	�-�1m��o�rrrrr}}}}}}}}}}vG�#ݑ�b��)�b��]����]����]����]����]����^�^�_K��bh��/ ^ �{��GA�R H�G@:c�1�c �x��G"�E�9L�Rն�KS�I��j|�>T�(lD�li����eF��i�i�6�M�#L�O�$j�$j�F� H�D@`��&q�Dd�(�kAUU����L��I�F쑻$nǛ���y�L`�c��G�#���z���y��`���R��R��r��r�M�4:q�m�$8�$8ލ�::�oI&��[���"5K"5M����s|F�ȉ�"&,��t#Tt#Tޑ��"c|'o�颪h�މ΄S��EkH�֑��#�GmyE�(�H�6����ԭ��!��B�D�',�d���X).�����6�aM�Sh+*)�)�V��+J�+J�-
�-
u�N9+G%8����Mb�LTa��1Q�&#Lx���;��wc���	ݎ�'v8N�'tK�Ջ�Ջ�j��R�T�mO$ͩRfԫ�Q��j]xڗ^6�׍�u���q\j8�6�VL��U��*�Ժ��.�5_�/◇qKø��e�&Y~I�_�%��	e��i}�_^%gg�Y��Vvx��g'�Y�j�5N)��F�
Ѫ��j��&���Ж�Z�kB[MhKi�	m5�-��'6���D��!�d�Z��j��)�+JnD���К���DJ851ZNrp��$�Tq�18�S�! ��mC�k�|�&٩��j9��I���,Ŵ,�,P"��F�B�|�p�?):u~NC�c�����+�L�X��8��!����'��1�ˤ�M.�S)��L@��mCq)�Ħ�7�X�Ji��SM��m���mĦ�7�X�Jmcq)��Ħ�me�Sk�նn$�q&�Lj�52�XcZ���6�Klc[c��6��X��ch;�N�Rm�6���ڦΣjl�6���Z�nk�Gk�j;^�QΎ5��[ָ
޵�V��y�M+Κq���q�[��k�K&���k�K&�h�iV�@��NV��8QZ���� �!:H^�p�+��b/x�ŏ�{J�ITC�I�Z|$���{��w������:��W��<�w��0�����A���U�$#x��"OC�H:�+]g��w��mxM�jK��x�և�R@`;|-8�Bo��:�j� �,�p>��b ��ľ)�\Mk���&��3��{�܉��L��7���k�I"�"�I�};�I��1������:�J&���m�	vH��������ܡ=L�������|���c�#�$G�H��v����|�>v����g������l��C[�-��+u��}�;1��l���[����j����a�� ���	��( ����� �� ���
ت�a�0H6؞��OPO �82o�sG�����h�!W4{�=��*�*�*�*�*�2�2�2�2�2�2�2�2�2�2�2�vG�#��1�S�3f��#0F`���3{9{9{9f�]��f�x���{Ǳ�{Ǳ�{Ǳ� ^ �xc0�b�E�9rZ��ն���9��
��(PaB�S�����R���i�M��&�i�� F��bi�� F��b�UH��čUCũ^�e��h��!�eG��� j�>@�����#v�l��F쑻L�7bI�L`��H�$}>�D��G�#���w�^F�I.X��7ç����"�JB6��v���jw�m^���!�y��x�Z<]�8׏%kH5�mx�C^6�tF�:#O7��ɡ�M����'B+^FƼ��y�����m�$�J-���#�����i��5*ȍ*���z�2tJm\w$��$��J�Ԍm�H,�ƽR��y&YJ�4�Fң+��dKB����S��w�k!�䢵�V��7�Z�+A�,4��ǁf�,����p���;��wc��xjAxڢ^6��f���jy|ڥ^�/R��i��b���mF+�Q��P��b��1Xm2�6�W6��ͩusj1|jG_��Ƥt��L�&w �;�p�^�%��Y���	�isx�\�g'�Y��VrF�хd�aY9Z5PV�T�U�5��&�V���Ж�Z۫Ba�И~�&�	��ctrLn�I���1�C)&JM�1�C&4�dƘD���͠�n9)6U���Y�hLP����#�rj���~iGɫm��Z���Zz���������@�I���LC�h�
��N�ݩ��|BC�c�W�WL-ޓ�+:`��.�&"�~,������s:����+<�YY�:���� :�ͱ�Vm�r�Xu�Zì��f���4����7KP�M-Cq)��1M�1�mCS��4@u�Z��Sm��Y�jefٴ[f�im�b�X��ch;�����F���5&ۃj�n�m�6���ڻ��Z�nk�Gk�j;^�QΎ5��[ָ
޵�V��y�M+Κq��d���ĥ#���w��5�ť%,ZRR�(�S��p��N!IA�Bt�����ɮ%,�����_�A�CBD�驓ǃ���������y�n�~#u���7x1��:���[�<�z��oP���#�Dn�{��w��k��:IFp����h^1+Q�i1�c�F�&���א���A�y�o���$�~Ӭ�Kk���mX����nZ�����?�S��#���Dh:-�����NP��u�j�7U9������6����҆̉��Sa�	��-�n�������P>}A�	��v�U��s�\����i������੏v�d5��L{�^헻t�����ݦ�~�@1��~����6���d% ����L0H'���������a��b�� )�-�D�)���ѐE�/�/�/�.��d{�=��)�b���#0F`���3f�]����]����1a�9��sGD � `, e��� 2�X ��9~Kr �ˠb!G��a�@c�t `, e�e�{.��t `,r�1��?`��G%�l*N@�9��
�'�(PaB�����R���(lD�li���lț�#L@�1&��2�����|����x�+��b���D0�����u�TCg��u�$nѭ�#vHݒ7ci���y�L`����G�#���x�@� L�&^��y��n�j$�R�R�9R�j%��N&��@\� ip>�� ����h����1e~�G;���.�w�sP�P���+^H��H��F�oH�M1���v���y��������F�F6��H��I5#f���4�5JA6�9B�����5)�y�F�;��)� N@��@�G+#d��]�S)8��ΣQ�����e�V<�+*%��l�`Q�"5���QZJ4�F��|���X�,�����o�'v?��p�ؼmQ/TI3SBM�<�mR�G��u�j]|֗^F+�Q���b�Ԏ�5#���ú:��.�mK��R��Ժ�Ԏ�5#��H�ø���L��Y{p�^�%��Y���	�b�+9<
�O��0���)��
k`�4�r�{���|[�ka�Ml-	mա-�J'&�ɋBa�И~�&�	��a������ct�RL���d"Rl��&�D����ۀ4��Bn��s�(]�&-	m5i5=hKi��MלD|J&4хd牥��i[x��&''Ye��Y�J��ǂ��=2�j�S+��DX%7N���I_�C�h����Y�%1t~+�����&�u�[��Vy����u��YX@u��c���e�q1/[��z�LK��bm����jf&������bm�b�P�Ƣ�M7h�����P�Jm�S+6͠��6�KlcZ��wkAݬmv��56�Q�6�T�pmSm��M�����spk\j;^�Q���׸�s�\oZ�+z�[֕�M4�:i��d5�lr�w���R��JR8֋���iIK��NV��8�$!I��z1�F8ǃ�����@�ֿ#A�����a�� �pn ����8]C��I��i7�M&��]7Z�F�t�k����	��7[�,�p^�14�]j@�(�!������@&�͸��3k���n�K|���O�:hmr5>$ݷ�iQ�ѵ���SzF�LޙX��?�9O�d�7_dm�DM�EIȌ�&� \n���9�M�Sa���Bm5F�h��WdF�k�����j�"?�ǻd5��U��s�\����i���O�X~
��n��@[�)�tǻe��{�A1�	��Ll��������da��ꀪ��a����'�19���Ol=�����ձT����`�l=�9��*��N�p�a�9�c��"�E������������#ݑ�b��)����3f��#0F`��K���K��b�v��: �!�C�9r�1�c�X�1��Xc�X�] C
=~Kr �ˠ ��9{.��tˠ � `,r��������90�ɆRն���9��
��(PaB�
P�(0��(lJ2�̡�(l�2�̡�(l�$g臊�	0<�j�$7h*8P��&q�De�De�Txl�&��>Fّ4�9b:ӣ[2F�m26� >�G�����`�y��=M�Sz��_�k��~կڵ�V�(D�(D�#\�T�T�T�#\�#\׏%5;��@	�GѪ�e�(�<Ф#A�$J֍�mD�]�K�s�ԻZH�����6��A�mSjH�ڍDm$cZ�����$�6��@�ڍDףW5�M�[�փ�4�m��6�ڒ.;��4�4]�#ȌD���0�=!=d�|�������Қ8䖎C&�%O�ˉE4KChb�U���+_k���������xo��w��[��_5�	�rL�ГmO8MIW����Qę�bM�GI�_�f���j��5^�/�e��e��b�1p��8LA�%��	e��Y{p�^�f N�'Ye��bv���&�7����isxS�T�a5AMP%��m�r[`��&�Aɭ�i-��'&>	g�Bq�(��%�����nC!�F���D.`�B��se�D���0Q�G�ct
B?:���L�T9%��s��">��q��Ĝ��M�A�MZ5P���Q<�hKn��͐�	��,���ρ�ڎBl�@�ȱ�ދhM`�
1�[Bf��|����U�) ���7�?�Ÿ|t����1�n�Z)!�$郂s�c��Ė�f�h5/[���:�.��5y�r�P��N��St��5�1�"�M^��7p15�9ezuZ��5j�M�jef��4��V��551Y�mq��k�v��:��b�wLr[��k�a�`c�چ�ww<�{lu6����6�P�?��1ݥ��q4�Q΍)d�7�zR5Õ;���q��N2�zoD��Z)a��:�Q��!|)睯	� �� 1��<T��d!����|u�e�,�t�-h���Nb�X�Q�����	�����z��u���T�j�Cih�\��,��QH��S7�eu�ڑ2։΂si#�m���R��z<ВF��'j���D�bD�$lH04�dI�l�Zr&���*lJ2�ĩ9մ]�-{a�	�i�ݪ�j�ګs�9����V����>>?{������tǻd�
�n�ۯ���Pl��/v�ݲ�i���Za���a��~����a��~���ꀪ�������;ؠ��U�{�=��sG�����h�4{�=��sG�����h�ї��}.���f����#0F`���3f��, e��� 2�X � `c��!�C�9r�1�c��!�C�9r�1�,r�1��[�[�X��G"�E�9r(�Qȣ�G"�Q�������=z�z�z�z�z`��&9KV�Z��ն' T��B�
P�(0�A��CbPٔ6e�CfPٔ6e�Cfn�*i����#Z���UH֪�Cv��ց"��e	@����5Q�bm��vFَ��:5�$n��$�$n���g��VսM�S{���7�ڵ�V�j��Z��_�o"�EH)ȑ,H�,H�,H�)ȑ)ȑ)�M*6��,��^B�W�s��B��^H��8ډ,��^B�K�sP�S��&ԁ��<x�<x�$���2Sw�)��^FN��5���R�hڦ���A�$\jTjTw\w hmIGP6��j$@�@��<��<��@��@��<��$�.�\Oy Wy1�R*o�Uͩt��˄�]�iVbD�4��ib��F���Y�N��k����Y�7���5\-��j\�548MI\&��3����bM�GI���3k�L���5^�/�e��e�&Y~p��8LA�& �g	e��Y{p�^�%������i}���&�7����Vrx��g'��=MPFT�� r[`��%��m�i-��%�_���91hN>%��cTrR7!��d# ���""-��pij�-Q���2��7m���h*nv��">nv��O-jd�1�5��MM�T�EM��:C)��#�"7��$&��"7���84�G��Ɂcu�5N!�`�g3$|87�b�@mƣ����D����4� ��zd�z������0�RG�cP�Jk��b^��P�Jb�j������|Oy��s�?�a�����c��0�Rt��9z�.�8<��0@c��!��X�&���Sm�ě:�.5Խm!S)���j�7�P��KӨ��Qͫ�)��:�K�)�6k[f�Y^���D��y��s�׏�K&���^��jl
׸�-�"޻���Pu5�p�NҒ�)���y�O���x���E ��|��A��V�Cφ�X�M\/!`��o����xrڅV�hM��5$�H>V/�;���
�M�M�b!żz�D�Z��6?�]cVÄ���&+DF
���v����V�I޸��h	,�<N���ɵF�����ȩ��ޒ(�GPp"_�H��F�o>�7bj5	b�n�L��I�6�M�(lKT%���
��B�
�`�D�*{��Z�v�ݪ�>s�;O�O�Z��>>>?{��گtǻt�
�l��_m��tPl��/v�ݦ�i����ꀪ�����������������������;ؠ���v9����h�4{�=��sG�����h�4{�=��sG��c�v>�`#0F`���^�A�3f��#0F`��`, e��� 2�X ��9r�1�c��!�C�9r�1�c��!�C�9r��-�,Q��G"�E�9r(�Qȣ�G"�Q�������=z�z�z�z�zn��w&�0�Ɇ	�0Na�sS�*PDT����¦�
�*l0��¦ġ�(l�2�̡�(l�2���>n�0P��X:|��ݡ�T:|����l�p�k@�kA��F�$jd��F�G[�6̍�$n��$�>@��$n��#i�����T�T�T�T�T�T�T�T�T�[�¿*��p"p"p"IRDWAE$EY�M*:47�
�Ck��DI�i���)�y)e�0��iy
5�k���j�R���K����(�� "Y !,�[����x�v�y)БQ�mQ�1 w$�H%bF�"I��iD5z�D�D�G�ǗǗ����wy� ���C�)�Nq�X�Y��8���M�����9��9��0�Ќ4�x�<H�%���w��1"1"1"4��1"u��:�)]gs�����ܻ���5
��8[P��3���j �5 ���& �g����i}�__������i}����'g�Y��VrxVхd�aY9VN)����ф�a5A5i��[ ��ʴ��V�۪�[u�K?|�ք��Q1�9)�JF�2��`�A�O8\���A� Pi@P���pii�O(jgb3�Du��yCh453���l"��ڙ<M����s���܍� �Q�ܒA!3L6u�""��Wn*a��O�J��t�RL�ګBs`rNl+JnO�ڿH�]�Q��B�|6���4+�B�]CNZ�` �>ki5�%~Eó�|���q���M�u�[a���'H~)rp�8�����91�mf�?�mL��1���D��$�h+&�AY�ɍr�Yk�ըjcWsp;�[A��1ɭ�S+m{X�.���7[��F�������SS\6����Qͣ�z�:�MCS1;�sh��޻��Z>%,���b�b�m�l���(D�!����ځk��WL��Ӭj/Q����^�?�A0v� �kE�9X^��� s���RŊ�u$���ֱ�'��F�p�Qܪ�!�γi=N0�Q4�.&�R�ީJI!@��!����N�L�$���|:��-a�R��Y�L��@��g���du�#i��g�� �n�Pؕ'���W#[��H��"l�P�@����	j�M��MBD�#r��H�JK\��Sw;U��v�]������������s�S�S�ǻt��{�^헻t�����6@1��0֘ka��~ca������p�p�p�p�p�p����������������˚=��sG�����h�4{�=��sG�����h�4{�v>�c�v3f�r�r�r��#0F`���3f�2VJ��X+%`d�����2VJ��X+%`d�����RV
J�IX)+%`������RV
J�s�s�sэ�IX)+%`������RV
J�IX�z�z�z1�1�1�]TcDcDcDcE��j��ܘn��u��s�`����↚4
h4�(i�P�@��̡�(l�2�̡�(l�-T��ܵ�>\@Z��ݠ��dt���TCf���5Q��F�Q����u�$n��#�� 6� ?�Ǐ�$�@I������ժ�ժ�ժ�ժ������������z����U�P�@��4wAE�'p	��u�$u �H�H��K��K��j�h�S�Թe�1�8׍�5����j�CǌOS%7�9-$��NYk^��{�����GkďHǘVa�+ƣ�h��='�Ry%�����đHHHǗ����
K�'����I~p��<Lw�!<����U�qNɗY����]S�)�V��գR��X򴬕�S8�)�%O-
m ��牤���]�b.�1#�O��g�d3����;��K �%�O�'����V{��уW$`��5rF\��W$`��S[F��Ʃ��T�r�z�j���>	���5��&��m�r[aZKn�Im�i-��'&>	ɏ�ra(��%�����`�DE�8\���<�"�)<MG		��!6�O"n�&�O":�mL�F���m��:�M����:�M��;r:?�ѯM�jf���O:��c��S#N�yA�W"1��b�E��̈́�iQ�܉7�H
"n���J�:��MŹ$m�1�`@u��Q����W-Ԥ����?��)�-MI&�����7kl?��mĤX>sc�m*W�.�0�ܵ�L��:�B�|�Eś�|�a�.,Ÿ�ۋp��4�Ř�-�m�j���15�cG�˹��צj�Z��)��sP��׏�f���Y^���G,����/Z��L7h��׸��v��54�9�6uZ���Q�N5��52�l��I����53�"tk��ծ:�Qc�t�Z��p;���e��A�����~�w��4�oC�
Ŵ)Q��a����G��X�Md�C@�L�ZUĳ���	�e�M>5��jC��m���*�(^G�9m$aS��D��D��y�x�� .[7����yz�P>`��y2<�L�ē$������둭�E
*N@MAqeqbM؛u�4
���Z���=�(D�$I�7)��M�Z�7s�]�WkU�|
|
|
|���S�������L{� �@Z`-0�ݲ�l�۠����4�Za�0�����l?1�����s�8U8U8U8U8U8Ulelelelelelelele�e�e�e�e�e�e�e�e�e�e�e�e�e�e�e�e���3f�r�r�r�r��#0F`���3e���2VJ��X+%`d���ǯǯǯǯǯǯǯǨ�������碒�RV#������h�h�h�����������������������h�h�h�U.�1�1�1�1�~�?s��Ϝ�|���&5S��NakaqkaqkaqkaqkM֚�4Zh4�P�aCM�64�P�aCM�64�n�j��T#����>\Dݑ�GO�:~�i���O�:~�je�n�[�F�m2<|���mV�X$�@���s��s��S��Sժ�ժ�ժ�ժ�ժ�ժ������z����U�P�A�'p	��"�"5�u�"*����Ȫr*H��"�)��!�Mi�h�V�m��F�oI7����EͩA�x��I)e�x��2jt mROgw���)�_�;�U��������"c�qIШ��\Kw�%���IB�"��5ı&G��0�@�Q��a%�Ǒr��aI�0��2Sz�)�R��H�w ś|e"ޜo�#iuq�R����+ FC�C-	`	D�ĢXbQ8Q(�1h5.�)�++V��+Jb�0ς����	ZV�+V��>
�o���9M�Z5vV�]��Wei-9ZKNV�Sդ��i5=ZMOV�Sդ���5��%�ք��Ж�%�$�sd�NL�����91hL?Zք��QH��Lj���R��B0��p��D�(�"5$F���[�����hF���#h+�6���vF�m�qS�`�֦F��� �ۏ
Q'�����u����)�X�h�ۏ���z�����$:�ă���u�����V ���+�� �:��c���4/-��:u���J��m\ښEޣ�����fc6�U�4�>^&���-:�!���|c�ע�r-/�J:��\p���Pu�ڿ�B�x�S-
�㨤�=2���'��լ1�M@�M��湸SmL� �N6�5(�sp)���M�Q�-r�YM����������jd��D��+Z�sp)��ֹG,���u�SM����rtwF� �K^�2�����f9,��sq�*"��*�A��$��	�N�!��2E�-��),����$�.۶�M�j�"p%�����'9�m�x�H�ta�y+��٬L.���2�j��0A~Z����5�q�N���E�jd�Dّ�bE���q���Z��0T$�D$��$�=S�>D�>hl�$�\@�\:�DT��j�I��j�2��M�(PaRr"մ\�90�:Z�0N�'K\��sك���`�j�O�O�O��~~���tǺcݺ�n��C[�0�L���l�cda�0֘d�l?1���UU�z�=m��[G����V�V�V�V� �1��-�Albcv.�b�v.�b�v.�b�v.�b�v.�b�v.�b�v.�b�v.�b�e���9r��-�,1�c��!�C�9r�2VJ��X+%`d�����������������������G<�9�� �ys�#�A��G<�Ɔh`ƆU.��ys�#�A��G<�9�� �ys�h`ƆU.�]T��Ɔh`Ɔhbc���~�?s�90�ɇ�s�kaqkaqkaqkaqkM֚�4Zh4�P�aCM�64�P�aCM�6	�P*lL�6���O��.#L@�2F�"nț�4�d�2�L��dm�fHݍ�H�<|��U��	5P7D�0\�-T�-T�-T�j��j��j��j��j��j��j��jަ�ym~Uy1�Et\wAE�T�$\�F��#�ȩ!;���(��I1�US��C���j���%�H�H���P:�ףQ5�oIYt#�\�JtsHae䔲�TV_�]����޿��r��5��bDV\5z������hᨒ"��"��"����H����-�d��.Np&$��!�	����PI���<ܩ���V�Dm~u��W�a5��NJ'=���c�pQ,2К�J%�%��`	D��X!�,��C&���c�[�䚜9&���d�r�(��9&'-	�Bb�М�Z�BsahNl-	ͅ�9�9&7G$����!��e$�I0"Bj�HMQ�	�9!5G$&�DnC��F�hDDZ�ʞp�PD����p�p'��F�i�hF�ErF�vma��vjf��l jf�F�l$�p3�� n&�ӭL��dӉ��.�~��tj�Z��2A� ��E���Jq�X�jK��Ԧ$1�d�d��M���)�����x���bi�$��qx�!�	����� o��ޅ�%aՠ�$�#���$§��uL��	��6�i��q�pX<���m��0��ʈ��W[���hS	53[��4���u�'�hF�6�ۉH9m��V�8'��9M�u[c�� � �"j�1z�	���>Q�-A�"LI��R�Уp+7�~hNOE7L8ڀ��!n�q�M�ʌ�ICRx���8_:C#��� �:?I'tm�(�@�AF��D%������-���Q"�mN}o������X�^G�&�2�>��,D��[���~n�~n��`�~`��T��P��D�xލL�&Q���dI��#v�L�O���F�P$l�m�i���ղ��M��"F�"$�FL7rcUmqkaqSfZӕ6%��&� n쁻��sw)����|�>v����cU���>>{a���0� 102&�6@1��OOOl�[�0�kd � ƘkL5������PPP[G�����h��z�=leleȽȽȻ��Ȼ��Ȼ��ػ��ػ��ػ��ػ��ػ��ػ��ػ��ػK�� 2��!�C�%�%�%�9r�1�c��!�C������������������A��G<�9�� �ys�#�A�1��]T��uTs�#�A��G<�9�� �y����.�]T����+��K��U.��s�\��+u��r�-�1:��0l�0l�0l�0l�0l�0l�0l�*l�(i����
l(i����
l*lJl*lL���t�SbD���"#�v&ى�bm��fDݎ�dm�NDӑ�c���d�����4�H}j�x��MT ����z�Pz�Pz�Pz�Pz�Pz�Pz�Pz����U�P�@��+���"���:H��#�GX�#���!;���#T�D�����	��M�
A;|:��u�A���5��Mz5Z6�Z@�������it*4������7���0�d��MI#�]��P4��3&�yrrI��.Mt��W�F���W��k�)XI-~x��8R	)���I�!���D�."t����M���o�ԭ����Xw�1x����a�9�Lv��B% @R )H������r����)'<���)1=�)'��$�)	@
BP���q`rBi�JM��I�9)6G%&������ct�RL���$#������#w�Dn�B�0��DZ��A�O8H��	<�"��D	�BDj9<u��Q\��+�6��ٌl 1��1��������y������H�nD�����5�7�4�6-��~�_��#�����@4/�x.+��Dx�>�C���hp���%��0�_��:���"71�w���tN���۽V��6�H�ܩ�F��Y�C5�?�Be��^Q'����'Г|�X���V����u#�I�0�rQKG-���e�oV�CI�ntNQ���|��Q�l_��q��D��M�f�W���
S,�2m���JMb�N�󩃐���A׊����@�B
LM)�K%�)�V���S,9��x&� ���v���@��M�tiZ�4?V�J`�$�$���D5Pmͯe%�#I��DKz�;�F����H��e� hkI6�G�V��Q�ui#��DU!U$[S�T�7n��ѭ8�'@�Wyj�ykB���պ�I��3���_�n��c������0`��H�<|�Cf`ӕ6%���O�'H#m�#[	� �s�;S�( `ؖ�%I��)�� n��pS�������v�m�T��6�|��T�l>{A0"L��d2��J�PP[[[OOOPPPl=���� �'�1=����NNNGb���=m��[G���������c�v9c�v9c�v9c�v>��3f��#0F`���3f��#0F`��`c��!�_�ߒߒ��9r�1�c��!�C���������h�h�h�h�h�h�h�h�h`Ɔh`Ɔh`Ɔh`Ɔ#�A�1���K��U.�e��Ze��Ze��Ze��Ze��Ze��N*�]J��t��uR��[�l;1��ƛ�74.H�+ll����hj���6��M���T�l�j�U6U�XZ�ake����XZ�ake���5T&9kM��e��}���[,>\F~�M�̡�*lJr��M�(iȚq6ĉ�#l�[�jd��#n�۱��4�@ ?�0I��ժ�ժ�ժ�ժ�ժ�ժ����0��X�*A�&��D��D��&�ȡ�g�y��QS��#�,GX�"��-��B�uȉ���H�H���)�����PkѨ��j�R�P���P����]�4��Yz��s�q�~�iz���J�#%g������Ў5I ))�A�K!E%��r��9$d��2LS�!)��%���hQ]4�WY���K��%Gf����;7��� u�c|L�~nVH�ŉ��4]�kE/� ��77�9<�BOy����D�9���"[:�Kj9	=G!'��%�����
8����3�.�:���l<�&���!���2t�Bn��M�I0�RL���q��">y�G�P�T
j�B�
84�
*y��8H�
O(�� ��5�D����"5�:���[��u�r�#h;���hS	6�0�hS	6�0��܁���S5�Z���?8�L�u�A�lm����$����8�A�x5��ԒW���l#oN���.`�OR���2�		�(�9]b�vR%��@�b;^})��N��h���2Ya-~���~)$�^H����[����ho��A��dt񤀸5b�ho��&��!�fڟ��S�s����N1��|�%������T"l%ȗ�V�Hwr����^��Jw�-0:�1?�� XͻqR���Pa��+�`x
S|�5���I7)"@���kcp���aS�����@ry�G�������6Jd��N_�,�LCr�����ܲ<���2Vw�o��i"洀�e�1dF��Bڏ6�%:*kѫ��j吚%�V�7�H�4�g� n���ւ���(U��~�6�F�Ěly5W<�����z�ě���m�L�7bnR%��t�Bn�*l0M�����r7*5::��$�E�h;[�������Ӧ�v�����~��n�� ��V��<&�G��=�|����	��&D������r��% �'Al5l5l5l<5<5<5<5@@@�{�ߘ�����'
�#�leleȽ�eȽȽȽȽȽ�eȻ��Ȼ��ػ��ػ���#0F`���3f��#0F`���3f�1�c��!�_�ߒ��=~K~K~K~K~K~K~K~K~=~=~=~=~=~=~=~=��������������������G<�Ɔh`ƆU.�]T�閆ha��ha��ha��ha��ha�S��R��]J�]T��uR��.ot�dj�i�4��ڥ%��
������%ڭэ���@�鋌�lϚs����>P�[><Z�\|��e��v���չ�{�7W&"(LDD�DF~�t�r5�����g�?D:~�t�bM�7X�>@t��i�4�e�j�m�����H��-A�Z�Ե#xV�7D�-T�*\�*\�0A�`�H�ĉS���r$O"�Ȫ�Y.p	Ԅh7���h�Cj@�ג1�$a�IQ�ISZH��:��uzF�h���&&�����I51����P���@��TwA� �I&�I���bTڒJn��%#�-�p��<o��)HK��^�M'8�G��襛j�OY)<��T���Ԓ:ͭr4)����%�9�d�OR
S&�)M�f��R�d�ܷi��Z�b�N]�:=��)��uG�N�a���7n$��S	(7�e��d�&�i�uG6`ku���&8I�?���&�DD�����p���?n ���>�O�A\��Li�DI�9��r"Ly����T�	��Ry�D|J!&<�#sLD��`RyA��F�JbG��D?8���6u��n���C�cz?�[�8��X,�&���۬C�q�Dj?i����Su����
è�s�s�D:�)$N�Ճj����a4�`ڴ�u��$�j#@��Y hmI6����j�Q�ͨ�漑�x�#��e�DDG�G�G�G�@�@���oT�Wy��M�d�<0��}&���G��oWb�8��O%����`OPWC�9��Nt9�+b&�@��[��T��&�؞�9�Nb%8"��	$�"X��I�o��ۄcC����:���Ԥ׋%3^ ��hS5��%tХ�Y<�޿,.D���c�QI��Rt4��N��c�Q-䨦�@��@�$����$�dI��"��#Q#Q&ԑs^�Dޑ�dD��N�*c|&�b&�bZ��nǓV�>�ϫ��S���y�S�@g��y��e�4h4� i�@�ae��6XH�P�(GT#���0�A��������`�*r���\���ϳ�S�S�S�L?LLLL{���=��10�tǺcݲ��l�D� ��)��Ll�cdS"������l?1�����ߘ�����'�1<5=����O~b{�ߘ�����'�A9���NGb��������Ȼ���eػ��ػ��ػK�����#0F`���3e����2�FX�`#,e���v��b'a���"}.�#,����RV
J�IX)+%`��G=G=G=G=G=G=G=G=��������.�]T��uR��K��U�2zd����'�OL��h�h�h�h�h�h�h�h�=2ze��Ze��Ze��Z�**TT��QR��EJ�]T��uR�a��w7���'��'��'9*[s\�i�n�˴�('n�˟&
l������?i��5Z
��鋏�ln���0�U��1=M��s��f4ܥ���M5E��ŭ4
�(��.>\Tӑ& �j�0<6�<:��M����b�$�۬(lʚr��M�"nѧ�5Q	*z�4=J�W�<|��v~�ɪ���\�?@������8�/��G�!B�uS���"E��A��y��6�΃h7��RSC��Bh��X�1d&�4:�4�A��	-xݭ a�yQ�Q�6�l,�.mF�iTiTj`�~���Mw���JC�%:���Q��0$�2Rt*!,R��IHJs�t�rs���yQLy)I�I 4) RH�Ԓ9�H��~&:��I������]d�:;)Z�%)����=����HmrW6�β��К�!((�%�.�ja$��n�es�n�	��L�`?���`�e������h'�[�<ݴ��A<ݸ���Ah�v(:ͅ9��G47aSqm�Z�rD�ͅ:�L�4m�h67�i�v*jm�h6	��6�lF���lr1ԫ���	���'�����
ly:��םL�H��"!�ixVH�HO'��m\F#�R&ŵ#h)���"k�0�QJ�$��k�R�Aܐ�ȩ��+"&,���"c|�\thk@ҝ��k��6GP5.;��,�.,�",�",�",�"1	.4��)��]���7����91~�Kz��D�I��"c�<��P���/Wҳ�ج�r)���'!��l��P���.����-���v�M.�'�c�1Y~�NS�/�WP]bz�6�Q⍍j�nbl^GQ�5Д�$�Yި.�?�ꉊr�5�@��xj�<Mt%����gz�K�q��dIȒq��;� wDm$a���h�y�6&���	ԅ,�$�Q8�<��_��ޙz�ާ�6��Ǫc��	&0y� l�m�l0m�����l0m�����#O�����i�4�ӐN@M9ն���ɆL0ra����n�>>>>>>>{a���tǺc�1��L ��L ��L ��L�02$�ȓ"l�cdS"���Ȧ6E1�����TTTS�S�S�S�S�S�S�S�S�S�S�؜���v'#�9�c+c[��v9c�v;c�v;c�v;c�v>�`#0F`���/ ^ �x#,e����2�FX�`#,e���v��b'��2�X�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z1�1�1�1�1�1�1�1�]T��uR��K��U.�d����'�OL��=2zq�q�q�q�q�q�q�q�d��閆ha��ha��hbTT��QR��EJ��	QK�auR��C#�߮�h��U'9�[vhr}T�����R۳C��'�M��'�����:{�%��M>`|�FP0��aST��Msan��\��\����OT�N\�rA=���T����G����|��U��֚M����ڭ������O�孅�
���>[�'O����t�b���CmS�mSć�����(6$�4=O��LD@~�3� ��<�U/�ѭ�ȩȉsȩ"5*�Ms|:К$T�bĎ�F��#��+"6�A��w��%
��C���Bĉ�";^@��hm@�Ѵ��Z6�j<���J֍�w\w\w\Kp),_�#Ȍ@h��$��CA5��o��K!�$�Q�a1�p�<���G':-x�
K��1��;�]N�R +��BJ@`3ơ�^G�C��v��4��=�@��ڕ��Ri������Vr��'PH������L�+�>	���I��Mc��n�m��S	&&���v*m���Z�I����~6���kF��kq5���1S5��.!��J@c�����qY���1�֍�h���6�[�F�k n&��"��	��H?$V-��w�5^8���pn\
#IRԲZ�)���ԉ�W��֟����Ԉ��}p7cnW�vމ�oD�,M�F��tl�
5�j���
v��(A�(A�op��!B��3-h��h�V��h��E�q�E�Œő�GrCl;� bTSz��˓W�	��rk����r%�\�oW2b�l��O)$��΅���ئ�s&��n3K����s%�S�i'#���� j�{)����f'��c��e~ �<�MI>�]�q#��3�q�ƢD
�V�s���Iq-�d����<RS��@�^G
n��7y⛼�M�x��h1	.;� ja܁�����ڍ��H�i#��GB)Њ�"bh���&&��&��,��,KQ8�<��w�@�"Mؓfݏ4�M�e���,i�j��F�ѩ�j}�F�H��i�$�t�m�l([aB�
�P��&90�ɆL7s��گ�j���������l>{a���tǺc�1��L ��n��C[��7_�n� �~A���u�Ȧ6E1�)��Ll�cdS�l?1@U@U8U8U8U8U8U8U8U8U8U8U8U8U9���NGbr;�V�V� �]�E��]����]����]����]����]����3f �x��g/g/g/g/g/g/g/g/g �����;D�] FX����������cDcDcDcDcDcDcDcDcC40cC40cC40cC40��uR��K��U.�]T���'�OL��=2zd��D�D�D�D�D�D�D�D���-2��-2��-2�Ĩ�QR��EJ��*$��\Ê�N*�/�g�NO�`�;=�v{D2� A��敲�1Al���j{������\��a����z�Ò
�4ܗ7S��7V�6�'=����sD�sD�vcaٍ�;u�~�����j�6Zۧ�ۧ�[��?s���l�"l; �
��NP{��'*>OD`���A�r#�+u��F�W�4% ?<6~��1q�#s��넌	�%��t�W	�S��S��Yo�̩�U$�PS�Q8�;�.5Cɒ%�5B�-T�F�S��_��$&�h���GkD�,��)��"5Mx�Si� �d&�4:��$J5I &)ݍ�m�F��
���gy�����G%�S@�K �"�s�1-~~ج��'��5��Mw����&��D�},�%YT�X�H.�=�Ԁ	�r��`5H�WY=�@�!JU���H�o@:�)���������*��� �T�ےF�W*n*a1i"<���mL�&�MGY��4�a1��:?��ڙ؍���ID&����1�dӈH�;��b3�Dc����l8R�汱���S��@-4�C�L�zm�z?7����zj#j�VA��D�{�1��Rt9��)�JS�iX �ݾhp5n��~�S�.YI�y�� �#V�-AdZ��2֎�R�[���7���EGB�B�BEGA65�H6���D���j��h��h���;��4�4]�	o$rs�Q1���{%�]���"s�Ȥ�N&8���s�l��s���n᫡�Ŀiy>�T�e7��1M���v')܉i'2�����}+:��'"r�l��s&)݄M�]H�5_�,�4���!��!�%:99�\��BX�&��W�J�V��ՠ��h4��,�"mI-h�#�����h��;k�my�65�H,�+ڐ��-����*c|T�HT���D�>AޙlǛ2�y�i��$��N6Ӎ����|�:F�#[�����nR7(��Mn&�[�9J��NR�)S���`��w9�����v�]�W�������s���	�	�	�t��n��@[�-���ke��~�E1�)��Ll�cdS"��G���4{M�G�������©©©©©©©©©©©©��NGbr;�V�V�\��Ȼ�����������������#0F`���3 ^ �x�������������������FX�]��>�A�� ��1���9�9�9�9�9�9�9�ƈƈƈƈƈƈƈƉuR��K��U.�]T��uR��K��U.�]T����'�OL��=2zd���ƉƉƉƉƉƉƉƉƉƉ�S��N*�U8��**TT��QR��D�TH\Ê�N*�K^ A�v ��'��� �S�Ob� }�m���eH�ob���@��h��(9.Os\���m�%M4�͇$�Ϫ��1����l	�.A��t�U�aه�蛩�&-���l�1�����5I�h�� ������U�U��*������칦扲��@lU�Z��MAQa����&���=M�uQu�b�u������F��F��y� �Őإ!";���R��*Hu+Ƞ󼵠u�7-v�&"y%_�j�$t.X��I4=Z�&]��I.t.n��/#v,J�ޠ
�'$��ŉjh�ƴl�^6�Yz�;�K�^���G"|��"hmH΄eȁ^���~�Y�7\��6��+�;�?)
�;۱&���5I !,��J@Au��I�},^�oR�� c��]�p.y�o�,���Hڧ��O�{Vi(������n�)<�&�ܒ53a!֦F���A�؍Nă��?Ѧ9�u���Lu��Ğ�7��c�4ZZ����?Z�Å� �܎�N'��H�ζ�~m��ML<�4�G���R�cZ�h_�!�q�.�sMYM	�[�'΄e�TC͈�|�B$ݼ��)�)�)�$�)�oJ��,�:�Be�F�I�F�V�0����"\�#T�D�*c|P��M�y�j#j5jH�ڍDm$cjH��@�bJSw�&���O���9�j$��Nw���D�{�9��M_��W�d������Sy>���
��D���5��bz�&��I·2r�l��r+<���'"��l��[!,���L�״�K'b��a�I)�x��mYޔ��8YTVw�)����"J��l�<��<��<��@��HƼv�����E:[�;z'oJ+"�ȩ�&�$թڷV�7���s�<��w��ݏ4��ڄm>@�O�T(�	#bF�"N����R�)C���P�(r�9��r�9k���Z�-v������sw;U��W�5_X|
|
|
~~~~~~~~�i���Z`-0֘kL5��*�*�*�*�*�*�*�*�GcM�4v4�ؠ��v(#�A��)�+c+c+c+c+c+c.h�4{�=��sG�����h�4{����ػL�L�L�L�L�L�L�L�L��3{9{9{9{9f�1�c7��������������������FX�]��2ǳ��"�###############%�K��U.�]T��uR��K��U.�]T��uR�OL��=2zd����'�''''''''''N*�U8�qT�TT��QR��EJ��	Q qs.a��8��UF%�`t
T	�s�:��>�4>�T b'��>�T�	WC#߆@�/ 2 U����#�A��'ք�M�G@x$t#��2�2��vrrl�.l; ��*�r~� "lT�1�e� e��C�/}.�a�'hO y@B�&��&��Ȝ�1�e@U����&4��7�d1�|�7OA�
�{�6P�\T�D6nq~D)�F�Pd�������&q�:)~F��Lh0[�C[�%����i��4��j��M�jݪ�-v�-���q5�5�l�X�#����F	G�t�SBH���`�b&�NP�HDp��},�ݜ���i��7:��Rĵ��F� N���/���Hܤkw���@\��[�kt�ڴƮ�剄$�O67��X���Sb��L�r4$�,Ί���:�lI`b�
w����&���-לDu�9�xq5�U�n��n��L$�T��Ź�%q�=�t1������wx��R�#�8R����#���Vn�Q�$<d�Y��:��;$�&�r��@��i���;u�#����Gꄛ2��N<ؼ�����C���N�P�6#�۽�В-<�j�X��Y*I��د�*B��#�ĵ9�kEH$���7���B�h���RA65�H5�lk��ב�ڍDڒ.;�4���˔�����ߌD��b�h�4�j$�<�i{)�_JoW����� �$�iw���ND�;�M��b~+�+;݊��c�#�#�ج�r),[t�L�tl�^@Ҥ�$#g��)�mQ��y�@��<Vz�6�0�@��Z���m�A�F��67�V���-��)��|[o�-�baX��&����}t]�t��~�A���w���L`�f@؍�F�#i�j�u>:�F�Q��4�tMnP�*s�9ʜ�Nr�9S���`�0v�;Lf�ك��j�Z�֫�����S�S������~~~~~~~��l�[�������l?[�UUUUUUUV�;h�i�����v(#�A��OO[[[[[[sG�����h�4{�=��sG��݋�ػL�L�L�L��9r��#��������������a���3 �,X�	`�%�K ��r�K��] FX�r��1�1�1�1�1�1�1�1�]T��uR��K��U.�]T��uR��K��U.�]T��uR��K��U.�d����'�OL��=2zq�q�q�q�q�q�q�q�q�q�qT��S��N*�EJ��**TT��Q �0��\Ë�yt��Ì1ዟ��
.��#�)r9���.��s(*EG/f�re,bYs�Fh����1�R ˁ?.)b�?c�
9~K~Kf ��d����T��{ٛٛ�{�v
h�h�h�h���@�O��ˠb'aJ�ߚߕ9
\�1b�f�2��[G�����������ko��֪��v£��['�OˣO�4�?s�9H�	z��l45\����d��-O@�Ac���~�L}�=�!�7�`T��Z�-s� �'� n�N@��b5��5�ꄍB�l1�P��<��T�?~�����9�#rTn*|2|�*}�;LM�J��PQ&�$�#�Z�Vp9�V)�BB�j��<��l���v����N'��'C�r֟D��Q��!��iP��9`Y7+�]��j{���C!	�3`��ۼ���u�/S��<��u�~�k�E��I�e�ޯ�\t:�����N--RF2��qH��|?����x�V��E�$ƣ���j�'	H���gr  i�zb�$�C͆��͆��͔C��������S��B6�D�>T$Ӻ���U@m���w�^�ۼ��0A�կϯ&��`����?�۴��Hշ�M��*A�(����ޔN�lkH�H�Q�ͨ�V�u+jFq�".b$S{)�=��ߍD���oƑ'�H�b����m� ��[,SɎ&��j w {;�=�H H ��^���#L��v%���.�	�4I�&�ҋZF���2taY�dj�G6�QD���)��h�ޔ[�;zQM[���±0�L+
��S�n��}t]�A�I�zc��f$Ӊ4����V�"��tj��F�ѩ���t�>F�#O�'J��R�iS���T�0v�>�f�pS���)�)�)�)�)�)�)�)�)�*c�1��n��@[�-���kt5��n�����a��~����a��~��������zx�x�x�x�x�x�x�x�x�x�x�x��������˚=��sG�����h�4{�=��sG�c�v;c�v>����K�	,X$�I`��%�������������9r�1��[�[�[�[�[�[�[�[�Xc�X � `,r��1�1��1��1��1���K��U.�]T��uR�WL��]2�et���+��K��U.�]T��uR�Ze��Ze��Ze��Ze��N*�U8�qT��S��UR��]J��u*�Uԫ�QR��EJ��**TH%D���8��0��4"�U.��eE�
.��0QtB��q�OED��xQtM�0��t��&OL��h�=G2�9v
.�P�D(b�PG2�9�9�40cDa���c0�ߎC�3{9 ����et�����~8�u����Q�_�@A�� ��Xc׳���rGD�v2�r}rvG�?S��4����7OJ|����}G�����t��!k�{Cu�a��[OLva�r��dM0Ll��/v�&6^�ձ��d5��1�f�0v\�~��]�϶�kt�~
�n�?.:�J�P0v\`칲*�`��1�L? ����R��J��a5��! ��A�4련b�t�u�j Vw����Mּ���`@�t4�
SI��L�S�VO�rC�ؿm
g�p;;�f�%�p=4�ݼ1������~u5���������Bm���M�p�k_;��J;8Bm2 F�4S�	'���\��ǔ l" i�&�(v�'�I����P�F�Q��4���@����ep�e��|��n�y�_���j�l^G�/���?��+��ݎ�v/ϫ�ˁ2�>����E�&�X�-c|[Y��
h���R�R&��h�т&��+j:(�@ �@�F���e�Tj9d�1d�1�y��6�j$iRI-�Ԋ$�{Z:(�6 �<�<�6	�{;�9���d�#e�"2t#.bz�k��,��׉�o�k#y���b};��1MN���#V�0���U4Z��U�0�L*v�NթϮ����?c�2�L��/��w�1��@���	tm>�?T�n�n�6Ӓ6(��5>�O�'H��i���ȓ�Kr�)C���P�-s��K]����i�)����~�?{������s�S�S�TǺcݺ�n��@[�-���kt5��n�����a��~����a��~��������zx�x�x�x�x�x�x�x�x�x�x�xˑ{�{�{�{�˰˰˰˰˰˰˰˰˰˰˰˱v;c�v>������K�	,X$�I`��%�����K �,[�[�[�[�[�[�[�[�[�[�[�[�[�[�Xc�X ��%��U.�]T��uR��K��U.�]T��uR��K��]2�et���+�WL��U.�]T��uR��K��ha��ha��ha��ha��U8�qT��S��N*�UJ��u*�Uԫ�WR��EJ��**TT��Q �0��\Ë��t⩖�<�Ĩ��@�C�0⩖�J�Q�B�����UJ��U*�UT��UR��UJ�q�e����%D0��@�C.a��2�-2��s�s�t����v�;EUUtcC*As�1tb(�Q���02�h�h�h�h�U� ����r���x#0�/h�aW����1<	��l��l>�PrOPv�9"?O<~�Р��le��m��� ��{�=m��[G�����h��zz==��OG���-���=��l#�o֛���l��C[!�������l�cdS"�l�A�e��M3(�c4����Ȧ7CS�s�S�V�+U�`�j��V�~
Z�l�_��	4�n�p�X��7{���9Jm��b��L�Lk��D��K��Ѳ�	=A�OWYHmZvy6����I�D��&��DH��u�q�H��:(�j�X�hQ5��j֒�u���:�j�_�PM
o��� &�$l* i�"rA��"{	�� 6���=��ȑ��78��uɃ�tj���5mD�����
�b<ӏ6#�8�f$݉6`i��v�n�闒e��p&RG���Nթڵ;V�7��PR1H`ŉ�Hn���|Z�4Tx�Pe�.֑6������Q�F�4v�����Q��Q��Q��Sj�GmQ����&�чB!�B!M���t3^:�ף@5䀚�G�ԁ��@��8��R1doYԆR�E�7�7�H�ELR1H[IRMZH��>���2�L�/#��2�L��.��;��L`M�M6	4�<�`�a�
�(F����5>H�P��1�A�@�:D�([aS���T�-s���]����ik����W���_X|���L?�Ǻc�1��L{�=����t��l�[/����)��Ll�cdS"�������l?[����l?1����zz=<e<e<e<e<e<e8�8�<e<eleȽ���-lele��sG�����h�4{�=��sG���� �1�7�7ӌ}8�ӌ}8�ӌ}8�I`��%�K�	-������������1�c��!�_�_�_�_�_�_�_�_�C%c�����覈����:�uR��K��U.�]T��uR��K��U.�]T���S(�QL��E2�e�)�S(�QL��\��1R e��Ze��Ze��Ze��ZqT��S��N*�U8��U*�Uԫ�WR��]J�qs.a��J����0�hEhEhEhE<��t⩖�<���ha��%]2���G8����2�ī�WR��EJ��u*�Uԫ�WN*�has�J�bTE� e��"8��K��@ʤ�A���K�K��UGUGUG]G]���G\�u�G]G]�12�T�����
�� _�_�C%`d� e��x������Lv~A�Oh���(>�O �l5���*��
�}D�М�#�b�[~A82	��sG���� �s��=lbc+c[[���yt�Sˠ�2�2�2�2�*�*��l?S�TS���ª�NGb��J�(T�2��eR�uJ�(D�1�;a�i��@[�)�)�'�)�tǻ`U�&��5Ap�܉:�i��N7@M��Iȓ]��HM�hI�*:�6��:	�&<���ᴘ]�%�+BN����6/'תe�M4�F�o'f��*ȵbI��b*���Z��ws$N��^MS.��§6 �-�O<Z���LF��H���95m�&�0��F�r`�\��[A��5mj}�O�(H#͈�b<؏6"M��f$ٽ[��v�n�闒e��p&RG���Nթڵ;V�0b�ޱ7�ϫ���F
���E[�2�B!My;^F�m#GkH�5�C�!�iv���^De�"2t8t8t8މ�����I�7��1Ќz: �{6�>���B!M�Qő���U�CꝫS�V&�!�"�F��X�X�j�G�����p�	�Be�ݯ�+��~ݯ۷�v�nޭ�ղ�e&��h6<�a{�@��D���S���5::����0uA�I҅�9J��NR�9k���Z�-v��LX�}a�)�)�)���0��tǻt���L{�@[�-��ke��~�_���dS"���Ȧ6E1���UUUUUUUT�zz=<e<e<e<e<e<e8�8�<e<eleȽ���-lele��sG�����h�4{�=��sG���� �1�7�7ӌ}8�ӌ}8�ӌ}8�I`��%�K�	-������������1�c��!�_�_�_�_�_�_�_�_�C%c�����覈����:�uR��K��U.�]T��uR��K��U.�]T���S(�QL��E2�e�)�S(�QL��\��1R e��Ze��Ze��Ze��ZqT��S��N*�U8��U*�Uԫ�WR��]J�qs.a��J����0�hEhEhEhE<��u*��S��Ze��Z�t⩖�<�s�ha�T��QR��D�TT��QR��EJ�qT�C�@bTC�.�e��W"J�UȎ4 eRZ\��˪�U.�]T��uR�]s�Q�Q�Q�Q�Q�_�_�C4C4C4C4@4@4@4C4@�4 �Ѐd����@`,r�{���;? ��dJ ��.s~�{/{/}G�
�? �]��%��c��a�-�D�1a�;D�1a��� �]��ˢs��tNc[.�lbe�-�AȻ� �14zr;�S�Vߘ�*�*���!LNGD䎉8b�ዔ�P2y@��+�̮r2�����<R	��l?1��l�[!���u��*��l��90�m�ﶨ)�����"lPJ��N@��l���K!��CT��HT\�ޘ)M#f����HkJ��瑭:`iS�y����dD\unD�t�I"[�9�h���PR4�Bj
� [/֫�#%G����769 D��NH����F��76#]��va#��h9��[@unF�F�Q��E	"��BH�l0y�lD�li��z�Pz�k����cɺǒe�~�A��}t\[���>��.��8�$��)ڪ���B���@��������M�GY�Y�Y�Ro�7��F�#v���u���!�:ȴRȡ�dP��	�o��7�om��Ƞb�����rH��#�8)#�:��F�I5Q8�A�גe�y&W��v�L��7{f�nޭ�ջl��@��ee�a�j� H��D�Hմ�h�ȓ�I�$�ri�� D���=S��ͅNl0ra�����v�]�W�5_X�}cT�l>{a�&&=���L ��l�cL5��i���Za�0֘ka��~�
�
���~ca����6 ��`R��(
�?S�S�S�S�S�S�V�V�V�V�V�V�V� �1�,N2ű�-�AlbE��r���]����]����]����]����2�2�2�2�]����]����r�r�r�r�r�r�r�r�`#�y��0�=�c�V=�c�V=�c�VJ��X+%b9�9�9�9�9�9�9�9褬G=G=G=���.�]T��uR��K��U.�]T��uR��K��U.�e�)�S(�QL��E2�e�)�S(��0��T��Hha��ha��ha��ha��U8�qT��S��N*�UJ��u*�Uԫ�WR��\Ë�qs��E<��<�cBhA�1*�Uԫ�WR��U2��-J��t��S��R��]J���J���J��**TT��L�0��%D0���ha�H%D�*�IW"2�*�2���.�]T��uR��K�au�.�����)S*`�L���03D3D3D3D1�c��ʘ)S�~h@2VJ��!�_�ߒ��/�}�g���l8������{�x0`A�K~h�=}.����a�9? �]��>�A����}.������ec(;A��FPr2������ec(9�D�11�9
c��9
�
�
�
c��9#�rGD�1s��́�
�'T�es�����q��i��NGb����LU�*�i��
���A0��qRr#w9����~
���6�r��T���H�j�Pw��PaP(ڂz5���l�-QzP�"T�#l�?s�;J�����Mݤm������մ
��6CZ��>}cM��>}@��c����Z�-v�;J�O��R'i��ڍvb5و�f9�:����I�$�5:�O�(I$
�a�͈�b$�`M�m6/�(/�5�f�l�M�<�.��:�#����n�����y7X�LA�~�NneNZ]HZ1HP��
YY#��E�&�V&�V&�V&�
F��#UR���$|В>2�>2�>2�j�S�X���L��B�E�B�Jss.��Bb�u����ݯ۵�v�n��~�Bb$���_�k��~ݯ�5�v�i�훽�iĚq�y�lG���y����	�H��D�#S�մ�h-��m�nQ5����m�Kl#N@M94�
��Z�7s��ڮ֫���>}�_X�}a����~~��L{� b`4�Za�0��������a���a��~�
�
�
���TTTTؠ��v(#�8U9��*�*�*�*�*�*�^�^�^�^�^�^�]�E؜e��X�1��-�AȻ�_R݋�ػ��ػ��ػK���F_F_F_F_K���K����^�^�^�^�^�^�^�A`#�y��0�<Ǵ�{JǴ�{JǴ�{J��X+%`d�G=G=G=G=G=G=G=G=�����##%�K��U.�]T��uR��K��U.�]T��uR��L��E2�e�)�S(�QL��E2�e��\������N*�U8�qT��S��N*�U8�qT��T��UR��]J��u*�UӋ�qs.bTT����A��cBhA�1�hbUS˭��R��hat��.�]<�ЊЊyt��UԨ�2�P@�E2�e�)���(碒�RV#��=<��"J���\�*�2��-.�]T��uR��K�au�.���0��T�Ɔ#�A��"�����������02� h@�״�{J�Ǡ��A���#��1���閛���Ko�s}f�r���tE��H蜅1��]��>�A����}.������ec(;A��FPr2������q�����]�csG�
c��9����h�4{�=��11�(\�]rr:%��9�A�b���2�2��OG���-���=��N~�鏨5]�0ra���逥�j��k��'�7@O�d�����H�WkU�D��C���$N;���V�-NDH�Gj���{�'�L{�CJ��5]�0r\n扲��-[T`乺��n��߭�����ȏ�0��|
|
�}a���M�L J�0�
�0��'�ݑ�"#s`����T�([a�����5:�N�S�
�a�͆	(0IA�m� �li��ݽ[��v�L��/V��lĚp6�����K��CU+ɪe$n]�`1bZ��*�0�72�j�I5N,Z�&�T�S�v���BH����<�L2�L2�?.�>�j����)��,L�F���W鋞M�N���Ӽ�w{Nٽ[(;��n�z�`m6�oV� m�M�m��b$Ӊ6"M��B@�$lI$�E	"��=�i�4�Ӑ"r@��'$ܥ�r�9S���T�$
�(r@��n�j�������������=��퉀����n��CZa�i�A����PNNl?[�UUT�zz==���v(#�A��PGb�;ض�[G�����h��z���ˑ{�{�{�{�v9c�v9c�v9b��� �1"�r���f�f�f�f��#0F`���3f��#0Fog/g/g/g/iX���iX����0�<�G��c�V=�c�V=�c�V=�`d�����2V#�A��G<�9�� �ys�
J���G<�Ɔh`ƆU.���0��\��]s�au�.���0��\��]s�au�2�e�)�S(�QL��E2�e�)�R�]s*@b�.a��8��0��\Ë�qs.a��8��0��\Ë�qU*�UT��WR��]J��t��\Ë��*)�'�a�ЃcBhA�Ң8��˭��N40�TH�UhbUS˭���R��ha�2�P@�E2�e����(碒�Q�:XƊTHD�TH%E8��L�0�C��U.�]T��uR�]s��\Ë�eR������.���MMMMMM��ʘS*`��^ҰX���Fo�.b��)�O�4�i��lhO �l5��^���W������9�A����K��]��>�A���Pv2������ec(9A��FPr2��TR��ec(;c�=��sG�����h�4{�=�bcOONNr[~b��ߘ�*��PPi��b��V��ثa��{�CS�L-[@��T��n���m�����Ɇ�r�9����sd5�	�%�᥮�=O�8����h(Nz�}�;.O?vD�{A���n�����d�Ϩ7@Zo��jc����$�1���?>}cU�����s�pR׹P&aP&>�D��C����9k���&�"[`��un�N�S�i����B<�P`���$؁���cջz�oV��lĚq&�I�i���\�n�w��_�y5L�˺˺˸�\S)#�)&��9�U9�U9�T��BH��$~y~�J�n�y7N:�8�����t�U�|1И���\�l��i��ӻ�w�b�cղ�ղ�ղ�ղ�M�M�M�m6	6"M��b<�P�(F��i�j��F�ѩ�j}�#O��Ȗ�D��76	��M͂nl0v���\�r�69��ͅNlj�Z�֫��O�S�tǹ�	�
`7C[����e��~���~ca�����h��z������z==�2�2�2���v(#�A��PGb�;ض�[G�����h��z���ˑ{�{�{�{�v9c�v9c�v9b��� �1"�r���f�f�f�f��#0F`���3f��#0F`�%�K � �����0�<�G��c�V=�c�V=�c�V=�`d�����2V#�A��G<�9�� �ys�
J���G<�Ɔh`ƆU.���0��\��]s�au�.���0��\��]s�au�2�e�)�S(�QL��E2�e�)�R�]s*@b�.a��8��0��\Ë�qs.a��8��0��\Ë�qU*�UT��WR��]J��t��\Ë��*)�'�a�ЃcBhA�..�US˧�N40a���<�Ɔ]hEhE<�q��O e���S(�QL��]2�et��Ɗ:X��G(�cO!<��A*)��8�qT�D��uR��Q�Q�Q�K��E<��S4 ]��ˑҪeQ��h`Ɔh`Ɔh`ƈ������eL��� @%�K ��r�����b�����dJ (=�O �82a�b�����L�%�<�Ԩ9�D�1�7��F`���3}3}3}3}3}3}3s3s3s3s3s3s3s8�3�s8�#(9b�����=m��[G����V�V�V�S�S�V�S�T Z`�l>�l>�N~�?TT�1V���*�~��[�ȓPl
�@J�#[�D�	�s�$MU���ʋS����fﲥ�M�S�*rh>~�@H��-�j��P~� �����#��4�S�[ (A@2���S����ʛ/���dT���505��l��_i��>}a�*c�0�������@�P��C��w9k���T�*r��H��:�[�-�ӣi��'0y9���%	(0I�i��lޭ�fى6"M��� �;�+����T��I�����Q����{Tb��������+��+ɺy���Lht7U:���K��U�L���e~�2�n�t&y#�������M������e{M�&��ӽ[6�V�'�Mզ���D�@IA�JP`��������t�:H�O���S����t�:D�"N�-�M�T�§6�K]��ك��Z�-v�9�0sD|
|
~
~
��L{�@[�)��n��C[/������V���PP[[[[G��������zp�p�ٚٚx�x�x�x�ytˠ�]�z�=m��[G����V�\���������������܋�Ȼ� �1��9`#����7�7�7�0F`���3f��#0F`��`#, �,X��@�=y��0�<�G��ұ�+ұ�+ұ�+%`d�������G<�9�� �ys�#�@RTH�G<�9�40cC40��u�.���0��\��]s�au�.���0��\��]s�a�2�P@�A( e���2�P@�D��$C.�rTT��QR��EJ��*)��8��0��\Ë�qs*�]J��u*�Uԫ�WR��\Ë�qs��E<��<�b��.A���8��C.�U2ys*�#�.�Ɔ]hEhE<�q���J��QR��E2�et����(碒�RV#��h�By%EJ��t��S���K��U.�]Ut��TS˩U0�BҮqP���4ha��ha��h`Ɔh�h���*�T���	`�%�����3}.�1Lr~Al2%�Ȗ�.[�82%��9
��3{9s���R��q�tN�9~h�3f�������雙���������������9�c�v9c�z���=Ƚ�eȽȽȽȽȽ�el�lelU<5��n�"l�.n��OOl�[����kd4��qjzSt�M׹��~q�Z�<n)�ͺ�0Oh0Oh*O\�v��ʓ�P8�2�0sh>{@��q�����w#�Fi�Ҧ���H���W���h9�_ZR�A*l�D��OG�T`���O3i���[���=��l�� ���c���}�=���s���)�)�)��X`�ƫ���7s��K\�NR�(���::�[��ѩ�jt�=�	�O�'Ĕ$��&���6� �7�vى6"M�M�m�����@mց$Î��/S��#���������.��C��пl�;�j��5OV�%�asհ�~�J�i�_�L��&^M������#�w��A�u�a�{MSզ���{M�V�͆	4�l�z�W=[���4@m��$��%'Ǔ����tm>:�"N��H����$�t�:D�"N��DܥNl-v��K]���ك��n쁻�h��O�O�S�v�t��i��C[�����PNPNN[[sG��������S�S���������S�S�S�Sˠ�]��-�AȽ�eȽ�eȽ�eȽ�e����������������Ȼ��lbc[��v9{K}3}3}3f��#0F`���3f��#,e��%�K � ����iX����1�+c�V=�c�V=�c�V=�c�VJ��X+%b9�� �ys�#�A��G<����� �ys�h`ƆhauR�]s�au�.���0��\��]s�au�.���0��\�(�QL���S( e�E2�QL���R�\���T�TT��QR��EJ��*)��8��0��\Ë�qs.bUԫ�WR��]J��u*���8��1**TS�O ��1�.A��b�q�0�D�e�g'&OFat��g)UO.�"�!J�yu**UL8��0ʤ�A**Uӊ�F40cC40cC�@ʤ�@��\Ĩ�QR��By��O!<���N*�ha��has�<�s�<��*��..y��WR��]2�1tb�:�;E�(�Q褷��`�#�E1�2' ���'?*N~T�)r��o�9
c�:'4tO�ǡ�@%��`�2���>�c�v>�c�v>�c�v;���݆]�_K܋�����O���� �11�9#�rGD䎉m�1�9�݋�ػL�������ӟ�� -0H7]�&9�LsT�{��1�	�0Ll�11ه�h��`��T�JT�h7ND��?s�(*?.�}�_i���i����7ra��ov�ݲ�n�ct/v�L<5<59���N~����������zz==�G��{a�2�2�2�G��{dU��i�� ��[/v�ݲ�n�ۯ��t0���v�]��sw9����~�>}�>ϟgϳw�k���&�"[at�>:��D�	4�l �@������āB$�`�M�M6	4�$�af$�ae���@e*��q��8�n�y&y&y&w�R��)]픯V��L�Msհ��h_�L�[�^�� m��m��m��M4�M4�m��m��M3�Vʠ6��6� 6�!���(0uA��$P�(G�#��b�l^�O��ē�q��ܩn&�*[��ʜ�NR�)����Z�-s�9J��NR�6>ρO�O�O�O�0��0��0��h7^�n���{A���L2
�l?1=����'
�#��S�\���.���]���L�L������������������ �1��-�A9r:$�tI�>��/}3^�f�����#7�0Fo�`��L�L���
c��>����9f��#0F`��� 2�X�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�Q��䷳��!�C�2�X � `, e���2�1�O�~8���%`���%D]T��uR��0��\�똎ys�#�A��G<�9�� �ys�#�A��G<�9�� 1*!�Q<�bTC.��ˆ%D0���.Ј���@�C�@ʤ��EJ��**TT��QO!<���O!<���O!<���R��EJ�qshe���Zhe���U2��L�d�Da�
.����4N4L��K.�d��E*��քUL�"�"�]<�yu*�\Ë��**TS��]s�`�HT��H\Ë�qs��EJ����\Ë�qs.a��8��0��S��Ze��Z\�� (ʤs���@�Uԫ�WL��]���Gh��E�=��r�r��d:��9�T�����������#�	`��^�Ac�t\��ъ�F*{9{9{9{9{9{9r�������˱˙{����#�G �_L�L�L݋�ػ��'?*[�lR�$tNcs����=9�����e�c���5Kb�b�b�b�b�oշ�����t�E�
�ӑ&;Zov�*c���~�Lv�_m�V�ݰ���l��m0Li�cLu  ��������s�9���Pi���Zb�1V��LU�*�G��{LU�*�~�_���a���i���[/v�ݲ
��??>v�\�W9����s�\�W;U�n�7s�����NR�)S��m�i�(0�A���	�O�'Ǔ�	Ѵ�"t�:6�O��Ѫj��F�Q�&�!%@m��6�@a���<�i�z��;�)]픮��W{e+զy��<�i�z��=[�^��/V闫t�d�d�d��M(�a�y��<�hl466� �l &��Rri�4�}�O�'ǔ#�4��|�:@�r��0��Z�-v���]��r�ik����`�0v�>�\���kU��W�5_X�}a��Ϩ>�|��c�1�� ��6@1���l�c`% �(A@2	��O~b��B��)�B�掉�b�v��v;b��� �1��-�Albc[��v9b��� �1�tI�蜑�>��3f��#0F`���3f��#0F`����
c��>��3{9f��#0F`�� 2�X�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r(��-�-�,1�c�� �1�c��!�C�9r����~8���������������������G<�9�� �ys�#�A��G<�9�� �ys�#�A��.y�.y�.y�.y�.y�.y-2��-8�qU**TT��QR��EJ����O!<���O!<���O!J��*)��8���2��C-�2��C*�TʦU2qT���.G8��C*�U2��-8�qU*��V�-U2ЊЊЊЊyt��TS��y	�)QR��E.���0��\��]s��E2�q	�%�0��\��]s�au�.��QL��E.���0��T��H?%T(��v�E�0�)�S(��F"�]GUGUGU��z(�Q��Xc7��GA�s�:�׳׳׳���QK�ʯʡ�/�?4 � �X�r�r�r�r�r�r���#�G �ݎ\�܋��_Rݎ]�]�\�����܋�Ȼ��Ȼ���ݎ]�]�]�݌�����©��P��u�su�se�e�e�L`��}�_f�ʄ�&H��ʛ	Mӕ����ƛݦ�i�� ��V���n��`-0�ݺ��u��4�Za���6��~ca�������{a����6��~ca����6��~b������a����6���L5��l?[�����n��=��0���j����4E�K�\�� n쁻���� n�k����iS���D��4�S���F�P@yA�'��=���5:�O�S���5>F�#O��H��i���i����������iD�iD�iD�iD�iD�iD�iD�i^��/V�6��6��&��&��&��&����i��P@�=���$Oa|�:Z�(N�'H������"tm>6� [��I�Lr`��f��>�X`�0}a���j�گv��������W�5_X�}cU��W�5_X�}cU����t��n���Za��i���Za���O~b{�ߘ�����o�9
c��9
c�=����9r:$�tI�蓑�'#�NGD�f�]�E��]�c[���� �f��#0F`���3}.���}.���}.���}.���f�2�)�B��2������������c��!�C���������������������������������%�%�%�9r�� 2���������G"�E�������h�h�h�h�h`Ɔh`Ɔh`Ɔ#�A��G<�9�� �ys�#�A��G<�9�� �ys�h`Ɔh`Ɔh`Ɔh`Ɔh`Ɔh`ƆU.�]T����8��0��\Ë�qs.a�'��By	�'��By	�'��B�*)��8��0��O!<���O!<��4 ƄЃ*�<�9���2�ī�WN*�U8��u*��V�-Z�B�B+B+B)�Ԩ�QO!<����QL��\��]s�au�.��QL��Bq	�S(�QL��E2�e�)�'�E2�e��\��(��G�T�u�2�]s�`�HE�������)�)�)���(�Q��Xc�X�]��>�c��>�c��K� ���K�ʡ�/�?4 � �X�e�tK��]��>�Aػ���bcv.�b�r/[O�x��܋�Ȼ��lbc[�r:'"�r.�"�r.�37373737"�!��zp�{� � ��s�9���[rG����������[���$MU���H���}�_m��u��l��A[ ��U����i���[�UUUT�zz=8e8e8e8e@U@U@U@U@U@U@U@U=��OG�
�
�
���~b����a��~�_����t���?>{cU����� n�U��W�5_X�}cU��W�>������C���&�"[arմ�k��������P@mA�	$���uB:�P��0�AQ�@�`��`��`�M(�M(�M(�z���D




̓�̓�͆����D

���P@�9"{	؍N�S����܉:P�-N�'J�I�$��tu:�O�S�q�&�0M͂nl*sDn
n
n
n
n
n
n
n
||||�{�^����s������~�?{�������kd5��l�����a��~���©«h��zx��1�S�1��sG���� �1��-�Albc[������܋�Ȼ��lbc[��#0F`���3f���K���K���K���K���=m�!Lvf�r���������1�c��!�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�_�ߒ��9r � `,~K~K~K~K~K~K~K~Kr������1�1�1�1�1�1�1��1��1���ys�#�A��G<�9�� �ys�#�A��G<�9�� ]T��uR��K��U.�1��1���K��U2�et��\Ë�qs.a��8��1**TT��QR��EJ�����QR��\Ë�qs.bTT��QR��EJ��*)�HD��HD�TS*�yp�ˌ�A**TS���**TT��QO!<���V�V�V�T��QN.a��<��(�QK�au�.���0R�*@R��1s�0b(�R�K�.���K�.���K��1b*:�:�:�cȟ�����뢕0R�E�����뢕0R�
h�����h�h��J��X+N1��N1��%�K �-�+@�L�]s��O��;#�=�c����������$�Incv.��7�7"����v'�Al�l�8�8�8�<e<e<e����������sd2��e͐˛!�4ߑ4ߑ4ߑ6C.n��n��L�0��da�l?[�UUU�c������$MU���ʚ�k���5V�9"Lvcd@5m�^�f��Pl#�b�1V�=@�@�@�@�@�<�<�8�8���8�ȽȽȽȽȽȽȽ����ȽȽȽlele=�~cdS"��������? �ȫu�~�>j�������l7{a����n��pSpR׹k����M�D�"v�����6��ڂ��$Ob5:�N�����i�4�|�>&�O������S��.F��F��F��$Ph$Ph"r@�m�!��éˑ�ꑩ�����P@�9{�6�N����@� P�����i�D��t�:P�"N�'H��I����u�#O�-��m�H9�0sD`�����0}a��X`���>������j���M�M�O�O�O�O�O�O�S S S S [�-��t��i�Zo�T�zz==�2�[G�����h�!�!�!�2�"�"�"�"�"�"�"�"�"�"�"�"��������v;��������������������ߐ[~A�e����v=��������9r�1���������������������������������c��!�C�2�X �ˠ����������������(����a��ч�Q�����Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�K��U.�]T��uR��Q�F4F4F4K��U.�]T��\Ë�qs.a��8��1**TT��QR��EJ��**TT��0��\�*�2���QR��EJ��**TS˧�O.�]J�e��.���<�����8�qs*�\Ê�0���˧�R��U8�e��Z�u*�uR�1��1���"~hA���*`�L���0��K�.���K�.�b(�ш���ꢕ0SE��Mu�uTu�uQJ��Ѐ�Q��똎���)S*`����������������c��״������C�4E*�4_�C��J��X � �%�K �,[���[��x#�Fn�.fnE�h��5���5�������zqzp�x�z=A���l
A����l�l�l�8e8e8e��kL5���l�cu��&���}����ݦ�P[G� [ -��ݦ�i�� ��U{a�i���Zb��z�{`e�2�P/P/O3O3O3O[G������V���+h��7!���!��zxʀ�u��ku��? ��>{@�퍑V����|�j����n
n��pSw���������^�r�Q7���̈́nq�$\�F�#r��H��Nr'8����P�(r�9J�R�)k���&�#s���\�:���&#V�F��:��j�մ	��� PT@��y��<���a�I�(G��6� N��Ĕ<؉(0y�P�(G�#i�$�t�:D�N��GS���jt�>&���r�h9.0rTn���S�"�4ENh���9�*sDT��������0}ak��������������������a�&�a�&�a�&7@[!���a��*�*�*��NNN[G�����C.C.E�E�E�E�E�E�E�E�c+c+c+c)��NGbx�� �sG�����h�4{�=��sG�����h�4{�=��^�)���-� �}/f�]����3f � `, e�g/g/g/g/g/g/g/g/g/g/g/g/g/g/g/g!�C�9 e���e�{.��[�[�[�[�[�[�[�X�1Fb���Q�����=GKGKG=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=G=��������������cDcDcDcD�C�@ʤ�@ʤ�@ʤ�@��\Ë�qs.a��8��1**TS��qs.a�HT��H\Ë�qs.a��8��0��%TĪ��S�a�S'��.�qT���T��N4L�0�閆=.y�iZ)Z'&OL��K.�],cDcDcDcE����2V8�#�8��V=�c�V = z������������~Uz�����ǯʯ��PǠ^Ұb(�Tu�uTuQMMM�����������������F`��%�K���~h�=~Kr��>�c�v>�c���v>��c����o�r�!T�T��(A��Ƙda��� � ����u�su����z����a���L24{M�G�_���e��~�_������M��L{��a�� *�7����AQj���;M�`���=q�z��E�
�T6
�	[!����'�l>{a�
`ku�~���������tS����Ȧ6��Ll?["��~�E1��i��["��~�E1��~A����'�|���5A `	�5^�W�U�n
T	�҇���&�M͂nȄ��&��76	��M̓�H�1��5m�C�'�l" Oa�m>6�$N��GS���E	"��=��P`�T:���'��=��( <���a�a��	6��=[*��օ�a�A��{es�����\�l��i�i���`M���V�~�A�ݻ�p6��؉4��
5B�P�T#i���}�$P��0�=z"��E�j��9*(Nh(O\P���=qBz���	�������s&90�mմV�(r@���$
�(r@���$
�0sD`�����#w5��k�����>}@�����P?��Ll�cd � ��4�T �����'�1=����O~b{�ߘ�����'�18U8U8U=����O~b�d �����'�1=����O~b{�ߘ��[G�����h��z�=m�2�)���-� �}/f�]����]����]�e�{.��tˠ�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�1�, e���e�{.�c��!�C�9r�1��{���x�1Fb���Q�Q�������������Q�Q�����������������������������������������������ߌ����9r�����ze��U eRU eRU eRU qs.a��8��0��\Ë����\Ë�eRU eR�T��HT��HT��HT��HhaƆhaƆ]2�0���h�U<���d��Y���%�˜�8��g��K.r\���1�c��Q�Q�E�3f���K����3f�r�r�r�r�r�r�r�r�r�r��z�1��	`�%�=~h�4_�/�Ǡ��F.�]GUGh���=z(�1�c7�����	i��N[~b��ߘ�*��s~���PР	���yA�*��VÙ�Ù� M
 �4(>�PР���	S`��V�Ce��e�Rc���&���T��	ǌ�'-OJZ���=)R�¥�	ǌ���*P8P�2P�2&�.&�@~ �������� >�*v_�;:��C��F�ȁ��n���jA&�i~�;�
�F!%1IHk��䴐��ָ��ɺ� Ow��F�-l.?s�AZ�֫�ݐ0sD`����$��7}Dn���	TPH���>{@����0���L>{@���?��L{��a�&=�~	�PH���>{a�)����j�A����d]��0}�� T��'$��F���95�Di���#N@�mrkh�ӐO\6������6��us����LT�LT�L\�L\�L\�n�z�Q�Q6Q;Ϗ;Ϗ;�һ�һ�ҁ�%w��w�y&4<��<��������WT󽲹��D�n�y�p%I�S��S�I4$��G��N�N��΄�΄�΄�	�<��y7X�l����z�d
	��B@ؐ6$
�a�m�#['�(O\Z���mQjڡ5Bj
��	�*PT&��MAP���&��Z��j�IȊ��'"*NDF���=Qz�4�Di�����#OTZ丵�qk���%�J��9*0rTZ��Z��`���Q���w5��ʏ����?}\�	`$M�J�ok�ok�ok�ok�ok�ok�ok�ok�ok�ok�ok�ߘ�����'�1@2
�l D� �=����O~b{�ߘ�����'�1m��[G�����h��z�=�e�S�"N���^�]��v���� �1 C��@�"{9{9{9{9{9{9{9{9{9{9{9{9{9{9{9{9r � `,{.��tˠ�] X � `, e��� /1�����������3r(�Qȣ�G"�E%`��GKGKGKGKGKGKGKGKGKGKGKGKGKGKGKGKr(�Qȣ�G"�E�9] ��~2��,r(�QȤ�2��*�2�*�2�*�2�*�8��0��\Ë�qs.a��8��0��\�*�2����"2�*�2�*�2�*�2�*�8�Í8�ÍNrG.r��9��R*9x��
�C1�� (c@P�?
�
�
�
�
�
� *(��e�d=�S��s���'��"[�8���J �46O7\��ݒ�O6\��7l?����[ a�����v��kdB`!3��B��6���R{�l�xM�`�&~�� j�@�Ǌ��23��Ȑ�tx��$&�$0P(L�O|��T�{#j���\Ț��U&�3%��sv�s����O��5[�.IS��[���W�ҥ��%6��Bq!R�郙�"3wb3pH��i��C�4����r���6�9��4�2���~F��"sz��=Dݝ�Nk�7%��HmA$6�� l,G�k暐I��n��۩�$�ВbhI1�l���ՑMd@�Y4ԃm�!z�m�� OR��	�B� �r�I=H�No^Mӻ|nM6�If��Kz&mX��������rz��$7&���AU9��l-[@�mմ\���Z丵�qk���%Ůj��;.0v\n������#wd
��9�(sTZ両�Qk��7&���BnMKj���'4-�O<F�8:�J:�2F�<&�xMAQ#M(���4�H֛At�Tc��Sȴb��~`\���P3� g�@�́�%?2|������y�~п?hy4<��<��U�#�N��U�#���C��Sպ����b�LT�*�(Gw�w�*yt4'W���M�Qq�*����~�jb}oD�� n�h�e��A��bn�$n�$�8�*Gk�^΃���E΃��.���M�GY	�X�%S��I48�8�/�,KL��/����`m��L�e���JN@�Ɇ�sw9Rr"��
�����|�j�M��I�' T��Bz"&¡���DÃg�H����"N\&�����$�9�P>P8D�2T�x��qRq�&��ն�ն�ն�ն�ն�ն�w#��G��mW6���CU͠��)��S�4��iS�&;Lv<��y1��c���cɎǚok�ok�ok�ok�ok�ok�ok�ok� � �(A@2
�P��dߘ�����'�1=����O~b{��1�S�1��sG��c�v;A�b���]��� 2�X�r�r�r�r�r�r�r�r�`#,e����2�FX � `, e��� 2�X�1�c��!�C�9fc#�#��)ؤ@�1��1���������������~2��,~2��,~2��,~2��,r(�Qȣ�G"�E�9GKGKGKGKGKGKGKGK~2���Ð���i�قc��M�1<'�/h�CJ(�@�ˌ�A*)�)QR��EJ��**TT��QR��EJ��**TT����By	�'��By	�-�����A=�{��Ys��W�t @��� �� d ?.  ˀ@0h`����C�{~��S��'9�l9%i��l�n��LP~�G(?{(?{(?{>D�}"j���������
��ρ����	����"��5��F�^�����z�[/Tke�l�Q��4����ys��A���Bq�4<ە��R�ԜwY)�@dI��
G��g�G�æ�EM׳��s�����g�����g��j����'46\�4��4ܗ7S�Q6�6\���6F�7v7i�j��(LNJ���19)�V�`����Rb9�L��y�{A�a)SdȚ`�4�$i�H���)D�)H�����7NDn���=qj���EM����ACL�U���&��Ϭ>}a���X~
T���=qRz���I늓�("*PDn�>N����%M�E������b�������"֚�6n�>s�]�WkU��v�]�WkU�|
|
~�?{��� SSLX`���� Z�S�"�4ENh��M�M�LX`���d]�-vA�|�-[@�=qRr"��DI��5AL�NR$�D�4D�4H���P`�T:����0uA��l0m���4 �(�Pl�ݩ�O$����p �7T�0hp�t5W<��SΆ�U��C�1S����nq�nq��<tڐ>��o����I��<�"ף@6����M�bz��@܍iA5��%�颠�h���l����/T���9�sIp�t5R�����鋞��OV� 6�!��"u��D�-2�j�s�NH��nr�9k����??>}���V�`�>}���]�V����~
~
~
~
|�j�Lf��W��
`t5�F�8`�1��n��=۠-7�t��n��@[�-0֘kL5��i��A@2
�P�p�p�p�p�p�p�p�p�{�ߘ�����'�1=����O~b{�ߘ�����'�1=����O~b{�ߘ�����'�1=����O~c��9
c��9����h���}.�a�;A��K�� 2�X ��^�^�^�^�^�^�^�A`#,e����2�FX� `, e��� 2�X � `, e��� 2�X �%�9G9f(��bXıG"�E�9r(�RV
J�G"�E�9r(�Qȣ�G"�E�9r(�Qȣ�t�t�t�t�t�t�t�t����XR�'��`��=�}~h{�Q�B�4<��B#�����R��EJ��**TT��QR��EJ��**TT��QO!<���O!<���ZZZZN%�(PO��G ���  @  �     2  1����������}{���^��ȓ��'��Os\�䩰���N<�N<�	�H(>�P}D�v\�v\�v\�sT�ln��O��
s�� �	�(>�l;44��6\����(>�N{D������.s~�`!�� �-n�$-N?N�2 �{��' \�rJ��x0`�\߮A�o��Vónh6���[[{����m�
�삃���q��zV���H'�Al�5��9��n��l�.l;1A��}�\�>NT�Oh?s@���f7_m��c���?sA��{���7�d�
�}�_g�H���9">rD|����#�$M7�M��{���7�M��i����j����v�|�Bn�j���V���n����s������~�?}����g���t��l��CZo֛���j�گv���������>>>j�گv�����|�*O\&�hPTT����`�?j�J��i�(0�A�J"Pa��D��%(0�A���	#MF�͔C͔C���	&"z�1�n�~~ǫv�n���<��<��/�:��%E�%CGǀۭ�㎃r�&���a䑹u�a�k�I��HT)HT(I����(~I�oH�ԅB�E�e�L�rw�:��������(4��>G�����[��Ӏm��M3�͆���C��`�L���4�4��$�A��J@�$P��0uA�I��	�*PT~
|�>}�>ڮ֫���7s�' Z��w9���1��L{���ݐ7vA��ƫ��0��0��10a������z�=8e8e8e8e8e8e�e�e�e�e�e�e�e�e����������������ȽȽȽȽȽȽȽȽ�S�1�S�1�S�1�S�1��sG�����h�4{�=�S�1��sG���c�v;A�b���]��� 2�X�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�1�c��!�C�9r � `, e��� 2�X1-�Q��1G"�Q���9r)+%`������RV
J�IX)+%`������RV#����������������=2zd����'�OL��=2z],�Y�Ԫ��U!8�qs��E<���ZJ��**TT��QR��EJ��**TT��QR��E<���O!<���O!hEhEhEhEvvT��J�(U���`Ӈ  1����~~�?_������������������}{���^�b����������.�.�)�lN{bs��؜���'�A<�� �ò��&�s�-�e�o��{��l	�h�� ��r��r ��3ng���
=.�]u�dSDb�d�E�@����A���*��vr[N{b�
s�<9����srsss~������@��	��h��\�1���*���[[[rrOl�_Pn�"n�ct/v�L��n�ctݑ�"?vD~�����#�dG�ț/v�ݺ	��Ln�cu��������4��?s���~�?s��[/�˵1�|�0PDT�DP�h(n�?r�����;e��}��[su���ܘn��w4F�h�����?L{�=����t��~�C[���j`j`	�	�����~|
|�ƫ���j�����jڣ���L{�=��Z�֫���P��4�ӐN@�=�ri�	� &���ri�4�|�:D�F�Q��j|�BH�$lH�y�lީ�l�@�F�ȝ���Nq�\�n�(F�.z�E9. n�5/ڧw���b9S�!��tk`�C��4Bkj��s�4̉�49 n��&*s8Z��H�6�~*r<Z��Z��`���q��#w�MPH5A �"Nhz�
_�E�N#V�#s���ܢkr�9����|�??(O\~
�l��90�9��*n�>}���@[!����kd5000��n��@[�+feI�W�i������S�eM1V��@U@U@U@U@U9��*�*�*�*�*�*�*�*�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�^�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�)�h�4{�=�e�e���A�b���]��� 2�X�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�r�1�c��!�C�9r�]��=�A�e�{.��tˠ�H�?.���@�*{G\ b$t�t�s�s�s�s�s�s�s�s�s�s�s�s�s�sэ�������'�OL��=2zd����s(8�'�UO.�]<�y���O!<�**TT��QR��EJ��**TT��QR��EJ��**TT��QO!<���O!<���ZZZZF�3hU2r	�s𩓗��@ d @ d @ d @ �A�3` ���0f;c�f9�A�`[ ��� �	r�%�`�-�\�	r�%�`�-�\(��a�)Q�!�%�֚4�8L��=��a��el�u8cel�{��0ȁ#��"� ^ �{�ː͗3�iS��-�\�{J�q82'!L[~A�S�1m�!W!W!T��'���59�
��r~����\�\߮o�7����T�!T��� ���������[~b�k�˲=�U����Ol=���Ƙ$lPOOPl=��	      ���ձU�U�T��s�<5<5@��l=�v�+a��l�V�퇹���Aj��F�ȏ��
��">[�;[/��
�i���h��~���#�dG�ȏݑ4�Z`-0�����l?TT[���a�~��[!���d5��l��C[�-��Ǻ`&=����U�zqz�=1�`乲�n��@S���ϴǺc�1��L{�=Ϟ��s���T����`�*#N��Ělz�*_��LT�O�>Ԃa�T:���T�`�=S��54�F�=�(?\�
D��5���mSu��E��eJm�C�	�E���n�6��~�>0i�6��7yQ�����7I#L#eGE���~:t_���뼍�w����6��F�n�L{hsh��9i�[T~�lPh#OT&���͍W��=���ȑ����m3/!75:5<�����By���I��j�V�'4'�PJZ��Z��Z��Z��Z�x����w#ɀ������Cg�M�7��7��T䭇�a��~����O~b{�ߘ�)��ߐ[~Am���ߐ[~Albc[���� �1��-�Albc[���� �1��-�A���#0F`���3f��#0F`���3f�sG��݆]�_K��3v���K��� `, e����������������������������������1�c��!�C�9r�� 2�X � `, e���@�*}~hvy��+����#�h�h�h`Ɔh`Ɔh`Ɔh`Ɔh`Ɔh`Ɔh`ƆU.�]T��uR��K��UJ��U*�UT��UR��J�����]<��T���Dy	�)QN.a��2�*�.Љ**TT��QR��EJ��**TT��QR��EJ����O!<���O!<��4 ƄЃ#Ȅ�ț`3  ������Ok�=�����Ok�=� * T �P�@
�}��L}��Ls�1Ls�1Lf�1����Ȥ�Ib��������D�	�8B�ڠ�c	�H�#� �RZ9����g����4K��h��/ z��1�K�A��\�s8��,�#0	`��_K��S�S�؜�*�*��[ ������=�				�)s��;A�dx"�a�4{�˰˚=���*��NNNNGb�ˑ{�z��r;�؜���v'#�leleȽȽȽA��d�4��6A*l�T�}hn�.O~bxjxjxjxjxjxjxkd�9P�d�`�ƪ�����?s@���f&;1��n�ۯ��+L��i���Za�0֘jz=8e8e8el�l�l���8e�e=��OG�
�
�
��������������UT�zz=��0shL�(s>}@��O���'����� ~�?{��������v�ݪ�-v��D��&��76-���%��ѭ�7W;��<�K�5N����k��h$�4���)�d��sJȁx�S?��#qQ�*0|��8��IO��X�>��⣎H`��g�h�-L
J:�j��JV��д��-6��4#��-A���_9�u���-53�ZjgP��Ρi��i��B�Sn�S:������x�S�N�C������H��Ǐ�#Zc[���(%([<`���q���yS�`����k����P	�!�W��WdG��>�|	U����%I�tǹ�&7A1���`$I��&D���	Sd���Cu����И�y1��z==��OG�����h��{�=��sG�����h�4{����������������r:$�tI�蓑�'#�NGD�����#0F`���3f��#0F`���3f���vv}/}/f��b�}.��� e��� 2ǳ���������������	`�%�K �,X����������!�C�9r�1�c�G/�X� " ]pc(�� )+��U.�]T��uR��K��U.�]T��uR��K��U.�]T��uR�O.�]<�yt����˧�O.�]hEhE<��T���Dqs.a��2�*�.Ј�B"����EJ��**TT��QR��EJ��**TT��QO!<���O!<���ZcBhA�0��q�w`IK��~\�r9xaH�
DR �0�A�")�{�{�{�{�{�x����3f,X�	na�;?.v~\�)$t#��1�c���R �b��%���U2� � `, e��� 2�X1T�9�4'=�P}.�v��,N��e G�	,DR(��������������9�R��	� ��1m����[~c�=�e����"�E���K��c�1�c�1�b'��e�g/g/g �_K݋���sG�������c��#�G/�o�n�؜��9�Rإ�H蜑�9�A�b����z���r�f�^�2��l\� ��`&�M��6 "l=�8e�~���`5leȽle�	��Ln�ct�����&7^�OOO~b{�ߘ�����'�1leȽȽȽ��������Ƚ�eȽ��2�)���r�37��37a�"�4z����L�����J�*>v<T�0��k�k��6�������"j�"-sTP�x��q���weF�k��;.0v\`戍<�y�4�ê	GT��4#[��í4DJ"PaakeqM�MAQRr#��U��g��ߛ��A�N��c@�����H�Ԛ��4�M_�C��8�Q�'�,5%Z^��	���+�Σ�Z^��8�6��ڐЯ���ޙ�=3�8zf8�?���<�8�C��`RQG��q�EG��q�E�HoM��0��1�r)\�nN��51l��a��sd��G�\���-�0N<Z�p�8�ʀ�`e�*�G�_�����PM���\�l�ce����ka��~��Za���ok�ok�ok��f[ �9
c�=m����"[~b�=m��[G�����h�4{�=��1a�;A�b�s�������������������� �1��-�Albcs��v>�c�v>�c�v>�c�v>�`#0F`���3f���˰˰˰��{�{���˰�� �]��� � `, e�g/g/g/g/g/g/g/g �%�K �,X�	o�o�o�o�o�o�o�o�o�o�o�o�o�o�o�o�e�K��h�����h�U.�]T��uR��0��\��]T��uR��K��U.�et���+�WL��]J�yuR��UJ��U*�UT��ur�UJ��Z-��0��\Ë�qs.a��8��QR��EJ��**TT��QR��EJ��**TT����By	�'��By	�-1�4 Ƅ��ZV��QC1� �=8zp����Ӈ�N�9.r],��t��(��`� 1c(�A�� X �  � �Q?@RV#��h�h�h�d�&W_� �1S��B����cȟ���뢕01�@�{2�1�OfQ=�D+ A��!M���ЂJ�lQ�$v��K��%�~h�2�FXUt2�#�a�!L[~A�S�_K�F]��@%�����2�X�]��9��v��t���3f�]����14{�=Ƚ���f��tN�>�@X$�ӌv2��tNC9�D�]��N0X$���37"�[�r;� ����sL��v9
br;�19�B�©ª -��G�M�ʓ*L����`a���u������dI��7^�l�b�M�r�����������������0�4� ��x�� �����:'b�v.�b�s�����'#�rGD����إ�b�-�\���9�Rs��v4ߑ4ߑ6 �2�^����M�˚oȔS�S�TZa�l�D� ��`&�M�� 6@"l�b`dI���\~q����D|����S�$M����|�ƫ��w#��"m�DM7��H'#�>[o��i�@�P���U�&PZ::F66H$6H$� ?n�9;(��GHޢe�OU��@�Q ���t�y���l�����=�s{ ���ۘ'�7`nonK`��E?-��}}0PP>>0j�5G��!�wB4�b@Z�(o��m��׺� �Ced�"5) �U��i�D�(;�D�Gu�M�y[�yeHڤ���4�o]�m뼍�I5�rF�NHmX���#R��z��OU��C|�#R=H�ȓ� 9��z��pd � �'A82$�Ȗߐ[~A�R�!K��.r��R�!K���'#�NGD���9r:$�tI��������L���L���L�K���K���K���K����3f��#0F`��K��e�d{�x"�����a�;A��K�� 2�X ��9{9r�r���1���	o�`ߒ��%�%���%���%���%���=z(�a�ч��F�U.�1��z�z1�]T����+�WL��E2�e�)��+�WL��]2�et���+�WL��]2�eu*�B*��˫�W.�]\��u��x��A*T�A���U�*�%TË�yu*+B)�*��E<����TS˩QO.�E<����TS˩QO.�BЊyB)�-���"� ƄЃa�T���Z'�R�K�`����U<���e,�ZV�B��Sʧ�O*�]<�yt���ʧ�O*�]<�yt�閆has�<�s�ha�T��N*�U8�qT��S��e���2�QL��E2�1R�yIQ
J�sэ�.���0��\��]Uuuu�� ǑJ��M��}.�xf����\߮A��7��<�c1��s��b�E�/ ^ �xc0�o� ��^�^�^�A�9�	-��'�Ȟ�"{Jǳ�������b�v.�b�}3}8�In�n�kc[����=�U�U�U����b�9�c�=��2�2�*�2� �9�
�D�	�dcU�����jzV��B�
�=A��
�$`��n����!�	�	�	�&�G� �
UO{T�r��y�-0uM	��ǟUT�>���������\����dM�3��)��fkc+b�'<�������b'4u��ǚof[�c����7�v�"��b��b��b��b��Cuء��P�vz���D�ޢg�Q3�����L��&~�?R����V e�q#�񻀁�� j�	��֫���d�F���jq"@4iA���M���Z�?7>(*j���#J�	
������BJq3�s�Ҁ6�t���xt��Pn@D� $*z�<��\�%"I�tI)��ZwmK%3id�ښ�%��Xjb%�
d�i0�&M"̮vQ,��R�&�|:�4c�"�Q�C���1�*9�nL
c55�V7� �Zc�͠�y�/��X�-A�n���[@�ru�M�Z�y�˭��^/��c�X�|:׏�Z�h�^-+�S�&9F8H`�;�q:�u��\k��'E��b�mT�Ӡy�@T�)s��o�9? �����O�9? �vG�#ݑ���d{�=��f�f�f�f�^�^�^�^�2�2�2�2�2�2�2�]����]��>�A����}.��t`#,e����2�FX���1���c7���a���/ ^ �x����2��,r(�1�:[�Z:[��9���9���9��B�����K����KG=.�1�d�cD��Ɖ�э'�Ze��Ze��Ze��Ze��Ze��ZqT��T��WN.a��8��0��\Ë�qs��EJ��**TT��QZZZZZZZZR�bULJ��U1*�%TĪ��S.�]<��t���˪�O.�]<��t���˪�ZW"�"�EhE\�Њ��r+B*�V�Uȭ��1�4 Ƅyt�C�@�C��hat��h8��˧�R��<���%UhET��UR��UJ��U*�UT��UR��UJ��U*�U8ЁƄ�Dd�#'�hA*�]J��U1*�%TĪ��S�bULJ�("2�#( e��E2�1R�yIX)+�F4F4N.a�Ȏ.Dqs.a��.���0��#�@1�A�"���01�OfQ'h[~A���rŰ9�_Q��"���_�@�.�� / ^ �xc0�o�/�/g/g/g/g ��%�K{J�Ǒ<���'��{9{9{9{9v.�b�v.��7�0In�n�nE��]�E�C.��d{�=�e��1LsGD�1��}2e����v9s3l?1��rT�Nl��9�i�A8U�e<�4G�J� �����M�:�Ő볼�Se�[/~=l�[�lb�[��'c�Xd'��-���AA���9�������ˠ�1e�)�xdi��������$��L@ѩ��M4���"�H�h!��q�<.5'[Rpյ'[Rpյ'[Rpյ)�R�L�S5
f��5�:�GBkjד[V��ڵ����mo�Mj��֬�Mz�~֬]�j��שޭz���"S���C��X��Պ�H�p: ޣ�BBN�07���z��/W����o�����6��Ԑ��$�oI��pn
��1ړ�hu��-��u<$7��r�_���|C��G�p'���:�m��y)�+�C���I7�tґВk�K�b�S���!'�ԁ�$H�$" ($(7"0""-##*(*F�������96[-�r�����Ó��eA�n|||�n�4�'�����ڃem9���r[l��4�ӛ����������a@���:`|HTnHTnHTn$FP�p�<���.r~A��'���r~A��'�����d{�=��vG�����������K�K�K�K݆]�_F_F_F_F_F_K�����}.��tK��]��>�@�2�FX�`#,e���1�c0�a���3f�x����/ ^ �����Qȣ�G(�h�h�h�����G<�9�� ],�Yt��e�˥�K.�d����'�OL��=2ze��Ze��Ze��Ze��Ze��Ze��N*�UJ��t��\Ë�qs.a��8��1**TT��QR��EJ����������*�%TĪ��S�bULJ��U1R��K��U.�]T��uR��K��U.�]T��ur*�Uȫ�W"�E\��r*�Uȫ�W"�E\���4 ƄЃ��<�Ë��Dd�]*!E�40���Ԫ�O d�	UZO.�]<�yt����˧�O.�]<�yt����˧�N4 q�'�<���GJ���R�bULJ��U1*�%TĪ��S�A*$�A*$�A**TT��L�0��`Ì.re,�D��\Ë�qs.a�R��K����J�IX)�)�+̢[~T�)��.��'��"}~���_�_�_�@��A� ���������Q��7���!�C�9{9{9{JǴ�����2V9r������e�e�d{�x#�G �_N1�����������"�d{��K��]�����!�������z��`% 1�1� ��$���1m���k�����7s����#���`�h���Ll�0}�_�fm�N~� "{=n��4��'���ߗS�'�1���� �2� ���������9#�9��}q�QG8a���_K�d�c*��.qq��˧�O.�]<��u**�V{U��g�Z�Pe+�\ʦU2��̮e�f��u���|�s yuq�B�F �(�c�@����:����¼%(�G�շI��r���5��ř��X)U���80'-�:E���gf�*A��A�"D�r� ��CCCCCCD�"ev�U��g�����U��k���V�U�B�d���.yq�HEsGD�)�B��)�B��)�B��)�h�4{�=��sG�����E��]�E��]����]����]����]����]����]����]���}.��tK��]��>�A�� ���2�FX�`#,e����3f�1�c0�`��/ ^ �x���X�e��E�9GKGKGKG=G=G=G=G<�9�� �y�e�˥�K.�],�Yt�'�OL��=2zd����-2��-2��-2��-2��-2��-8�qT�Uԫ�0��\Ë�qs.a��8��QR��EJ��**TT����������U1*�%TĪ��S�bULJ���U.�]T��uR��K��U.�]T��uR��K��W"�E\��r*�Uȫ�W"�E\��r*�Uȭ1�4 Ƅq��ҢG2�ʢ�Q<�t��̪8��˧�R��<���%UhE<�yt����˧�O.�]<�yt����˧�O.�]8ЁƄ�Dd�#'�hA*�]J��U1*�%TĪ��S�bULJ���J���QR��]J�qT�C��K.r\��YƉ�S��qs.a�S���K��UG=����SDSD2V=�A�R�a�>�c�=���ȝ�0��<1x����/e� e��o����������%�%�9r�1������VJ��X+%`c��!���^��F_Q� ��K��9�	,X#�F`��������`#0FX��/^d1����f䎉�bc-�J��\���֘&6*N�s��%DM���e�۱#M7��|�<�ܚ��s"Dj$M���ާ�πTZo֫���%�����=+d5��rT���[2�*�쉰�y0v����T�����e�".��8�%eV��̮es*�\ʭs*�ZTT��Q �	Q �	Q y
� �r�U.�]<�yu*裍*qQ��G�*h\�$H�"T�䨗\�s�@*`e�
\��c�����k�ē�U����é�����������u�.a)x�+]K��"�_(�����7��O�����UBeu*��U�1�r�	K�2]���K�!hEh]<�<�к�
�'yt��UR�QJ��B+�WQ�E*c�B�" �pc*��".Ј�B"��\0��QJ��-N"�d�*�<��]� �sG�����h�4{�=��sG�����h�4{�=Ȼ��Ȼ��ػ��ػ��ػ����K���K���K�����}.��tK��]��>�@�2�FX�`#,e���1�c0�a���3f�x����/ ^ �����Qȣ�G(�h�h�h�����G<�9�� ],�Yt��e�˥�K.�d����'�OL��=2ze��Ze��Ze��Ze��Ze��Ze��N*�UJ��t��\Ë�qs.a��8��1**TT��QR��EJ����������*�%TĪ��S�bULJ��U1R��K��U.�]T��uR��K��U.�]T��ur*�Uȫ�W"�E\��r*�Uȫ�W"�E\���4 ƄЃ40�TB��
.�0��'�2y�Qha��˩UL�@����"�]<�yt����˧�O.�]<�yt����˧�O.�T��HhD]�v�FU qs��\Ë�qs.a��8��0��%EJ��**TT��WR��h�h�=.�],���Ӎ��UR��U8�qT�D�D��9裑G#F�9] C=�`���v~A�2'g�#ߎE%���Kr��-��e��؎]���(�Q�:Z:X������2VJ��X+%`cȅ%`d�r�1�c0�o�/�/� �����K����iX�r�r�f�f�r�r�`#�2�F`�����%��D�]��V��;c��u����*�{�]�(A�e�b	���R��
'zr���bޔ%	,Zi2��4��B�'��b�+]�zb�7*�u�uA��4BG���4CU��Ё8m���F��{���>���}G�������ж]�Db�uS-2���e���S(�QR��]<��u*��Ԫ�WR��]2�et��S(�QL��EJ���A�̮eS-R�<��O2��Z�v�U��h�E�� G�#�<�)ٽM���Q(�?N���a���mĘED�F7�'��`�H��k2��fWu8�k�ļX,�dD�b�4=�T]���]8����\�s9�={9vsG�
������"���G@: ߎC�/{9{9{9{9r����,~2�G"�E�9r(��1��懲�#���A����u�	]� �11�9�A�bcs���� �11�9�A�bcs�����Ȼ��Ȼ��ػ��ػ��ػK���K���K���K���K���K���K����3f��#0F`���3f�1�c0�a���/ ^ �x��ߌ����9r�������z�z�z�z�ys�#�A��˥�K.�],�Yt��fOL��=2zd����'�Ze��Ze��Ze��Ze��Ze��ZqT��T��WN.a��8��0��\Ë�qs��EJ��**TT��QZZZZZZZZR�bULJ��U1*�%TĪ��S.�]T��uR��K��U.�]T��uR��K��W"�E\��r*�Uȫ�W"�E\��r*�Uȫ�ZcBhA�1*�t��h]�a���U*�Ɔ]<��T���A*�B)��˧�O.�]<�yt����˧�O.�]<�yt��HT�v�E�hDeR1*)��8��0��\Ë�qs.bTT��QR��]J��u*�UӍ'�OL��=8�J��U*�UT��N*�h�h�UG=r(�a���G!���] X�{�9�D����?�K��r ��?%�U~2�r�G.�r�r(�-,RV
J��X+%`c��X+%D)* �X+�9f��e�e�dx#7��I`���"{JǴ�{9{9{3{9{9e����K��]��.h�aQG��h�Kߚ)�9�����P~�AO��5V�(
�h���=���JD�[��d�a�M�D�}H��Ui=~�%�^p1ʙH�'����Ұ��Z:)|p]�E$�x5d�mI�֫���
c�ni5����k�A^E�	��Sߩ�֫����@$�uԨU!TʦN"�E2�et�����e�_�ߎ_�ߎ_�ߒߒߒ�4E�h�h�h�h�T��G8����U2��� C;D�1 ʠ^�_K��)Rs�U TO{.�11��9��A��sF�S�ۭ6�'7@��ܴ�����a��:ړ�hc������۬ͻn�H�\)ZL�hQ)�M!�ТiI2;p�����u��
ʄ�`
�������Zi�i������M<�A�����R���	�H��(%"O8&�qA����K[(����&���&�A�`�c���5M�e͗�M״�h6@1����%J��4'�\���8����.PР	�8�1L[�=�S��
h�#�rGD䎉��:'$tNH蜑�9�A�bcs���� �11�-�Albc[���� �11�;c�v>�c�v>�c�v>�c�v>�c�v>�c�v>�c�v>�c�v3f��#0F`���3f�1�c0�a���/ ^ �x����c�
9r(�---������G<�9���K.�],�Yt��e�̞�=2zd����'�OL�0�C�0�C�0�C�0�C�0�C�0��S��WR��\Ë�qs.a��8��0��%EJ��**TT��QR��"�"�"�"�"�"�"�"�TĪ��S�bULJ��U1*�*]T��uR��K��U.�]T��uR��K��U.�E\��r*�Uȫ�W"�E\��r*�Uȫ�W"� ƄЃa�S)b�.1p�(%h�.�.�=<�yU+D�Y����S˧�O.�]<�yt����˧�O.�]<�yt����-2���.y�2�Ê�WN*�U8�qT��S��O.�]<�yt����˧�O.�UJ�q���U*��Ԫ�U0��S��N*�U.��z)+%`ƈƈ���� e��_�@��c�dNA���2�^e��)�h��K~2�r�G.�r�r(�-,1�c��!�C�3r�2V<�2VJ��!�^�^�_K����������$�I`��qԨ>�����������c��;A��cr��T��b�嶆�����͡0Ȕ�'�l� >.H�p��-8̩�ޔ%5��z���F��}_L$�0)�~��H4"Wy[�9L�m����V�F��8\I�S$��! *�b.<HBҸ�8�	m�jV5?,O��&��y�u��Gsa����\� -�1��c�C�; hr ����B���0J�A*s���y1�Rc���5I�Ǔ�6]�6]���?[2~�\�l���s����H��H�Go�[/�Oݎ5]��*r2T����)B�R4�q��#��6����l�8m��@n��-Ot6DM���Ht��:D6Z&B%��+�Q"8���?�[��"���F�*��kW,�i4���m�&�B��"o
�$�nhQ4���`lX5�&�����}2Z�\M<����c��e�I��$�N$Ovs~- p������%��I�kj��*sDn�?}�V�-PTZ���ɇ��w&�"j�ϝ����i����~�?n�ۯ��&6AZ`-0���״���L�V�S��b�c+o�-� �����o�-� �����h�4{�=��sG�����c[���� �11�9�A�b���]����]����]����]����]����]����]����]����3f��#0Fa���3f�1�c0�`��/ ^ �x���X�e��E�9GKGKGKG=G=G=G=G<�9�� �y�e�˥�K.�],�Yt�'�OL��=2zd����-2��-2��-2��-2��-2��-8�qT�Uԫ�0��\Ë�qs.a��8��QR��EJ��**TT����������U1*�%TĪ��S�bULJ���U.�]T��uR��K��U.�]T��uR��K��W"�E\��r*�Uȫ�W"�E\��r*�Uȭ1�4 Ƅкe-�!C8ĭH��N�U<���e,�ZV�B���˧�O.�]<�yt����˧�O.�]<�yt�閆has�<�s�ha�T��N*�U8�qT��S���O.�]<�yt����˧�O.�U8�Í%U<�yu*�%TÊ�N*�U8�qT��9褬��#"�C@�?��/}�0-�A���*�*�*����h���g/�����X�^(�Q�9���c0�a�����3{3f�r�������������e�e�e�������#�Ԩ>�A��L�K�K������܋�Ȼ�T[��kM�
@|\MmU�$�2�OTP
�7.�-.�#t �#6���kT4�BS .�4�8��������~��������ۺ��d�)�M c�վՆ��L���~Mx|�:�7�|����5��u*��6,E��5�x���ı�e`Yy�r�]N~�-�>�\M<���	�Oհ'�NOh��(j��>N.~�q19+e=+u9���Q���%�K��5V�5\�5\�'j�0N<�N<�NJ�NJ�NJ�NJ`�d�l�jq�4�$jѪI�G�eě#��΃pN�pN�pOS��4���mױ����`!$�a#�������"2E1=�F<@���qx+[���;,׊�L�p���*E�H>KWؼ;�CA	j�6$�CU3�J�X�������u�S�y����t0u�~~��?Pw�S�����D1D�r��kt�L�Bz�մ��ϳ�i����n�7s�>��Z�֫���7s�9L��l-[cU�|�>v���[�v�ݰ&�2$T�����=��2�l����ŷ�ߐ[~Am���ߐ[~A��sG�����h�4{�=lbc[���� �11�9�Aػ����K���K���K���K���K���K���K��#0F`���3f�1�c0�a���3f�x����/ ^ �����Qȣ�G(�h�h�h�����G<�9�� ],�Yt��e�˥�K.�d����'�OL��=2ze��Ze��Ze��Ze��Ze��Ze��N*�UJ��t��\Ë�qs.a��8��1**TT��QR��EJ����������*�%TĪ��S�bULJ��U1R��K��U.�]T��uR��K��U.�]T��ur*�Uȫ�W"�E\��r*�Uȫ�W"�E\���4 ƄЃO*�K.q��\��h�Eh]J�2�e-+E�uR+B��Z\�� e��WZ�U8�qT��S��N*�]8�2zd���Ӎ���R��U8�2z],�XĨ��@ʤ�@ʤ�@ʤ�@ʤJ�eR0�he*$.av�FU qs��].�1���2��qp"럏Q�C%cٔ@�1��4tKa�'��O�@	��lrsO{a���ų��{9v~A�d1���a�G�/^�����;
�f�^�2e�e�������/���z��=m����T�q� ���^�f���2������7d�T��z�{��xɃ��ja��Đ��������eȩ�#~I._�m�9����N')ܞI���5�Bp9$[Uae9�il�	mU���'�[A\�����<��n]�L�?,C��N�m[���ۯ����$^A��,C��b��KΥo����W�kH�LW6�a�����'�	$�kGI��m�d��[(r@�9Sa+�˱x��b��t��)�ͦ|�О��>ODD�<&��y�0��~q��*O\`���r"D�v�+u�<Z�D�.F�0��\���	`〡�NPI�du�zas�5m�"vI��ܞMP���g�S��q�5�$jaS����iR۱���V_4����F#���u7������»r���B ��H��PiI"L+7%fԞ"+��3aؘ�X��#Q��vn�� z�C:
�H�̖�%w�V�$Mש��U̍�(����[\HZ�F|)<�@�kL㼡��JP���J<`��?8T���n�*��-O@�A�s��J�S�����l�Ϝ�W+t@5��n�ǋ^�Z���4o����邁�!��zp�{� �����'
�
�
�
�
�
�
�
�
�������������h�4{��9
c�=�e�d{ٛٛ�v>�c�v>�c�v>�c�v>�`#0F`���3f����=�c��=�c��=�c��=�`����/ ^ �{�?c�?`��G(�h�h�����G<�9�� ],�Yt��e�˥�K.�d����'�OL��=2ze��Ze��Ze��Ze��ZqT��S��N*�U8�qs.a��8��0��\Ë�qs.a��8��0��\Ë�yt����˧�O.�]<�yt����˧�O.�]<��uR��K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��r*�Uȫ�W"�E\�ЃcBhA���N�8��e,��V��SʩZ&R̥�=<�кy⩖�J�bTFZqT�*Uԫ�N*�U8�qT�D�D����%�̥�h�=J���q�p���s��c0��S��N.a�S��qs!8��U qr#�1����2����0��U.�]TcC�K��Jǳ(����9q � ��F]��A��������扲䉰���*��1م��T7A1����C/e�`O��3�\��a�A�o�1�1�4{�=�Um�������Z�\�v��m�:c��nD�\|�j�y�L}���"[/Nj�*-[T�l
���*[T`�0<���#l �*.���5�o�W,��,�)�
5	�5�P��=d�k6�)��ő���	еn׶��i1��)��PiCp'����!�vn$i�ܽZ��x�Y�^��Ќ����f9�xZmă��H>mޯ��z��W�~ۺ���ZY��J���+��c��xi�'v�:BK�ԍx��Y܀�$��#}y7s� �?<�������� L�$?.�?8H�T|n
H�TD��wiS���*NA��*O\~�j����'� j���%-r\T���8$~0m�pm��6�hz�l�"r@MmSȴ��=�T��7�-sY6^F�OV��#`e�@H�i��iݤn*8�����za�����|W����yG��\�Q�F�Z�H�4��Ь4��rbD�Nmͅ#ZD��+�ƫ�3�#+��b�$� ϟ������3�c���̑6��܆��#L	�>P<&|��sANH��( H�e�J$`��(&�hP~��"7[�'�-l.>v�9��>s����r�>ۮ��ku��{���[/�'������9�A�\�-��?Sߘ�� ��'���1<5=�����OO~b{���c+c+c.h�4{�=��)�B��vG���/^���K���K���K���K��#0F`���3f��c�1�c�1�c�1�c�0x����/ ^ ���������Qȣ�t�t�s�s�s�s�s�#�A��.�],�Yt��e�˥�K2zd����'�OL��=2��-2��-2��-2��-8�qT��S��N*�U8��0��\Ë�qs.a��8��0��\Ë�qs.a��<�yt����˧�O.�]<�yt����˧�O.�]T��uR��K��U.�]T��uR��K��U.�]T��uR��K��U.�]\��r*�Uȫ�W"�EhA�1�4 �ʩZ'L��K8z��yU�t�V���)gR�R�N4L��Kq�0�Y�Ӎ��UR��U8�8�8�8�z�r(�Q���Fh�c̪�h�h�KGKG9r(�a�ƈƈƈƆh�h`Ɔ].��y��2�q	u��s�#��4 �z�z���z��)T�;D,1�#7c(3sG������=ۮh5T4��?r��KS�"i�"i�0[A��O}vOl�.l; �i�ۮV땦�l��/�˵��n���ŹBbG��Zr���V�7�	�j��T�`O؍?T6~]���"i� j�-O�-Ě���ϒ��0����>D��m@��RE�W�Ad���.�G+��]�B���sxYsu�����nނ&=UO�Y���O�p���7Q����P���P��C�r�J�m��:6�`PiB���n&���֍Mhצ܍�-� pk�0�L�[��RQTp�h+����R��:D�8�����4��%b���'<�B"rHݽsS��6�(�DO&�u��fԑ=���5mF¥��S�S���v0}��ߊ���M���S�(l.LJZ���L �t�B����é�F�̒&?2�7Gj���**Nh"l$L�Nw�-����I	��� �V����l�m4��c��?��~��8u��0E��������ւ����V�"�J�u��4��ּR�ƳB�`�I�
���Լq/��ʔ�צ��"@i���8j OS��I��^E!4�6��5b�F�w��?.�{z��*O\�n�0r\6~(H��l�QL��d��4���q�p�U�T�O&;0�=�d�u���?s�_i�v�ݺ�M���Ovr��[8��7 �[Pl=���l=���POOOOOOOOONNNNrrrrrrs~�
�
���Q��їїїїїїїїїїїїїїїї��{Ǳ�{Ǳ�{Ǳ�{����/ ^ �x��,~2��,~2�G"�Q�����Q�Q�Q�Q� �ys�#�@�Yt��e�˥�K.�],���'�OL��=2zd��C�0�C�0�C�0�C�0��S��N*�U8�qT��\Ë�qs.a��8��0��\Ë�qs.a��8��0����˧�O.�]<�yt����˧�O.�]<�yuR��K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��ur*�Uȫ�W"�E\���4 ƄЃ�=8zp���V�V��Sʧ�R�N�K2�e,�XÌf0�˱��`�4��Z''L��K.�\�Q��xa�1��00�?�3.z1,bZ9ȣ7������^�^�e��X�e��X�e��X]U�RV
J��.�1����1�, e�e�{�F`���^�ܟ�N ���2�)���-�18l�5�5�
~��ku����SeSbTؑ6Pn�n�#l Z���*{�@4��`���=u�j�t���1qu�u�M�7XF����%M9!��:y�:�$T���F�5H�r���$hY	y.7D�{-s� ��S��j�|���dFeHDq�`�y�z�T�K��#���☔$�h!=Q��m�B��x$�z��:
x�ׅ7g	5��RP^V֦��#���D�%��1d�Bn��M�I0"Bj�JF����Pc��A<�G���!�܎� ��h47aq6jdi֦F��a�L6c����HqR�A��u�)&�kR(�d�֥kޛHY:�gC�k�婥��W		���ԥ���X^�3HB%�6�B�r�jYF�6WH�[�чf�L�6	$n�xhY7'rE���1d�~�J�><F�>J&�O�%"P`�T��T`���8�|���m1�m1�x�Ț����U�C�S�Ry�3��ūf	��֘��s��<H�m�~�i�<�Tt`D��yޙ֣��p��>�f8t�C�գ���:�#��\���D�r���WW�'¹�V��*�sx���D���F:�����'�7�HM�I� jȈ�ސ>d���Ԑ%��:��6@�n��yA�+���!%@m���S�C�iꑭ��i��*NDH�e�Zy���s�'�l�j��g����">v��"j���?s�6��P}cumSeɡ��=١��qA��� �S�Zo����f6_Pi��u�a��l=� ���`��l=��S�Sߘ���Űշ�-��
�?\߮o�7밫�����=��vG�#ݑ���d{������������������=�c��=�c��=�c��=�`����/ ^ �{�?c�?`��G(�h�h�����G<�9�� ],�Yt��e�˥�K.�d����'�OL��=2ze��Ze��Ze��Ze��ZqT��S��N*�U8�qs.a��8��0��\Ë�qs.a��8��0��\Ë�yt����˧�O.�]<�yt����˧�O.�]<��uR��K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��r*�Uȫ�W"�E\�ЃcBhA��˙�98�q-)�Sԧ�OR��=8�d乘��G���
�CG/G.�C(b�0�锲�%�F������1�^ߘ��Ƿ�=�0 �dz9���E��!��@
��1�`s ��� �0Ȝ�"f �:c��,�GA�e�U����A��*�*�[i�.n�44� �{�]�&9�n�"l���}�=�S��3��f���� F��5�������m�[(�[���iSa�M�Bm��l"n����ٺ��u���<`�"� ʑ5cg�#
��x���#���,F�,��)�I#X�"�GPY._�΄ �9Bu�Py��#\�"Dց�R.M#O7��"&7�lmG���D�%��Y4��%��R��	\j�4�F�eaK�J;��	�Lsp��:�nJ�saZKN%�ք�Q1�9&7He#��H܆B0��ΣA�*!��1\�5�[�\�G���`�h;����l1��֦l$jga�vn��vw��9�vpA�V�X�6�4���8qG�+j+�gf��vo���rv:���H���A�L�5#Z��'z�Բ:hR/	��)���uQ�u"��&��N�a'�Ԍ1܁�j�Ow�Q��m }X�_��5�m��f��RH���bF� P�ˉ&y�:
�I(�m����5D��Fː�um4HT6�r>�`�MoMA�hzm��8����jC��FjN0�Y�m-I�zc��!��jJգ�x�w�Ŵ<^ WZLr�i�*WZ�J�_7��Z@��Q�+WZ@�kx-\CA�Jjk�`~�ST���'��u�A�I�ε*�_��d4���	N"�ЭS�!4ر>'�&���.�j�������W����"����M�����(�[(9J��m6(0�:T��j���J��)H�g��k��S��fS� ��l;.l�%s~���n�S�&-���e��}�m7�M��}�ݭ7�M��}��m��a��{ca����T��'��?\�\߮a�A�@.A�A�®��d{�=��vG�#�F_F_F_F_F_F_F_F^�1�c�1�c�1�c�1�c �/ ^ �x��ߌ��������9GKGKG=G=G=G=G<�9�� �y�e�˥�K.�],�Yt�'�OL��=2zd����-2��-2��-2��-2�Ê�N*�U8�qT��S��qs.a��8��0��\Ë�qs.a��8��0��\�˧�O.�]<�yt����˧�O.�]<�yt����K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��uR��ȫ�W"�E\��r*�V�ЃcB~�b���ĳ�fNL��KJz���Y����)�����C(c��)�����c�:�" ���2�Ok�ߘ3@"} ��O���dxdxW�� ����@ ��9��d��NvA9��dI�ȁ
��\� ����c/��� շ�{�h�nh�X��[l;0�=�����mrb����
���ӐL[cu��[�S孖��F��?a!���@ ?����#i��I�4����$>�5PjǍ�X�H��-�ʯ"�����~UyW�9�$yH:���9d�A�QIN�R�"�7����z��$k�����"&�m�h����6��$��<���j�TSy")�f��"֥X)VK���t��L�)�S~�E/�)U�sβ��a8���V{x��+F�ςk�����'6$������^p�Q(��!��%#q�0����AQ�h0y�G���&���s@��h:�gQ��m��6�Lc��qn]��y�N������8I�uޯMf�&��h;)ښ;m�|+�Υ2ɴOh�SnN�� bV����"�ܬ�sb����C�`tQ��~�4�Je���W�⚔�~�ʒd�7�I�I(�Kn�X��PI(7��Ԙ��OI7��ҙ !�q�D��T�׉���y�5�S��3Z<|t7X���[w���W	VJsS��YI,�����"�1�oL���D`��p������1���+��c+F3x�7�"Jo�uH�o�5�r�4R*cB�`ܿ�JgZ�ЮY��pi���)�j$��hjbǦ�ъQi³7L��m � �Su�B�68��-�j�55�0rl�F�qXS:ԭ{RV�`�@]$�I(�� jɲ������^NE5��|De$`��s��O	&""O�9��I֫����Ol �9"P{�9O>[hl�� ~���z#��Ӑn�Zn����l��.v˝��l��.v˝��i�cL`�����(>�A��A�A�@.@+ou����9�®��d{�=��vG�#ݑ���d{�=��vG�#��1�c�1�c�1�c�1�c �/ ^ �x��ߌ��������9GKGKG=G=G=G=G<�9�� �y�e�˥�K.�],�Yt�'�OL��=2zd����-2��-2��-2��-2�Ê�N*�U8�qT��S��qs.a��8��0��\Ë�qs.a��8��0��\�˧�O.�]<�yt����˧�O.�]<�yt����K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��uR��ȫ�W"�E\��r*�V�ЃcB �3�q�32rd乘��8�q-)�S�'(�~� f�@A������o�g��^ߘ2�9�T��М�9�+�^��h��Ps��@ ��{~���wg�No�9�\��=��ݰ�l-�H6�l9 �rA�8<	��[ ��f-�A<	େf7S�LOD|���9˝��n���k�-��5S�Z�\T�DZ�@�=F
�Zh4�&�avD�$>�H����dH��7�0��F�d�=L5cg���7�č��Զ�(��"�N�E��$J����SD��E� �E��"� �4F��O;�����X��Y�R�dIoF�x�4;mF�bTVw�4�P&����JEB%=L� �,�H6�R-�Q���5�F8M'���K�ʧYY+�j���u��8LO�° r��0j�5N%������~�&>	������,�hL?%�	D��D�󈏂!s\��-�J�p�������r0(�uG	(�� (HyG	�BBA��h+�ۉ�x86;ۉ�y� ���N�΂4yG+��c�����M�M53c�""1����o���1��I&���mԃ�r�1����R=7h�"1��֥M=5��@�)�kV�
ܩ�$�y֥M+�Z:�#���F�i���DJ	$��ԑ��+7��"sպ����U�4ԓ+�V��Gu��Ʀ�*�p~:��"�"Wq<TKG��G^$ �V��;<[�ѼH�'��X�+��D�n-"�r�7�� �:�.%��L�'�R����BQ�I��j+��q�nR'?��h
��P�q��qFC�,u6�p��RD��Q�(��ǜ��k �D��� @rO:�M�(п1�	��j׭MMU�ft>�V�f�QD�A5��m"T�%��[�ɴxS|De�ގ�P�;Q�:��Z�7v�4�5]�7�U�n�0PD`���A��#t���v���~�?r��Oܧ�S�)�����˳.�l�1���ó�l;1�5�5��
�
��N}������)�b��)�b��)�b��)���d{�=��vG�#ݑ�c�1�c�1�c�1�c�1���/ ^ �x���X�e��X�e��E��������������A��G<�t��e�˥�K.�],�Y��'�OL��=2zd��閆ha��ha��ha��ha�S��N*�U8�qT���8��0��\Ë�qs.a��8��0��\Ë�qs.a��˧�O.�]<�yt����˧�O.�]<�yt���K��U.�]T��uR��K��U.�]T��uR��K��U.�]T��uR��Uȫ�W"�E\��r+BhA�1�{J 3@�tE�̜�9]��2rq-)�S�'(� ����J�@ �� * U���0K�c���9>�[vhOrJ��q��e���	�o�';"NvD����&9����ow L[}b��	��'��OsD��Pr���+a��s��:x+aٍ74�'����>��扦�n�O�0l�0l�>P@���s�9KZh6Q�O���7P0l0���֚M��M�DM�Bm�4�M:4�H} >��۱��x��7�L�F�.�tO"�OSx��I�_�]�W�U�Ut\u��h$��I �#h:�M#R����-����j�ELy΃fSDMѲ�i-H��>���A$�DmHGk�&Ѻh�Sw���DRy0���SrמnN����Iu�d�Ht\�mR�IUͪ�	��м,�I��ed�����S�Ҏ�,�p��8LA�f I2�����1'8LI�{��|�+6ɭ�QH�MPxVք���">%���&�(�����%#q�H܆B*!���q�P�&���O84��B��v���J�Ğ�y�E�$��wCS6��D���?���ؿ:��GQ<H�+�N���D�6�����I�[�G�@�禰RƇxp�X�3���㊕dC�<�� �Ĳ1���f��-�lS��{��6:��~5�γc��;8Ƣ����m!1ZW;��:�<(���J^�A��kP��(�����܁~�Ԥù�Q���\W(�����ۭΥԐ!��¹Dy�-���� +�ČY�Ն��+��Ar�nv4+
��a���R��i5�;x�Qơ#AL��R"�qx+��1��},�����xXX��c&��P �֣����f�n*`b���:�cS5�դưX5�3r.$�-I�SJ�H޷*pN���S4�L�.8Z֤�,�BDn�Kd&!��k�$6��$��m!4���jF�%�]Ap5!R�Z<bPp��Z�$lQ�:5�F��M����:�r�9ګv���n~�?r�V�ջun��l���l;1���Ý��l;1�5�5�m��N}���m�7똦9
c��9�c��9�c��;
�
�
�
�
�
�
�G��c��=�c��=�c��=�c�� / ^ �x���c�?c� 2��!�_�ߒߒߏQ�Q�Q� �ys�<�s�<�s�K.�],�Yt�'�R̥�=z0�cDcD�閆ha��ha��ha��U8�qT��S��N*�\Ë�qs.a��8��0��\Ë�qs.a��8��0��]<�yt����˧�O.�]<�yt����˧�O.�]T��uR��K��U.�]T��uR��K��U.�]T��uR��K��U.�E\��r*�Uȫ�W"� ƄЃc���@�  ����H??"{����aH�`�3)e�Q��?.���s��''dNNȖ��-��[s\��=�{�$�4I�h���'��OsD�sD���A�x$� ����T�T�T�T�T��'�S�X���d�l����l��n����i�[.v땺�?s�9">rD|䉪������9�r#t�F�ȍӑ�"-O@�=�'0�>Z�*l0���CM6�!6�!6�M��(6P"l�D�au�	��b:Ӓ7ci�����@?�Ϙ�>�ڵ��~[IRDWA�'p	�ELS�1N`��m�QI\���NUX���DO"�e$Fd�����k����m��΂+���"���dnS����,nT�Y�Ȓ'F��J�6�H������r��\�kQ+��J浊�m\m��ۨ��a�s��hV6�]F���R:��)�ڌV��Ơ�������,�$�NnK�����)�:�nO���j�����4`զ�&�+I���rc����&��GÒTrBj�
MU�I��&��C�a��!���"�F����.�Q�D�84�G�A�@Ph�p'�[�=�� j9<IG4<� �<l"h$�ǂ$�4�� y��o9]��AC�
O_����4;ۀHy��s��W:�Ca.�n��p	<�%"BQ,�"L*����i�jJָp������P�:�7�sJjB�@pW����&�i�d0+py��$��W���jC��-�u5'´qx�ۈ:0�������R�Ԉc�~�u�5�r�R���u�ۓF�bx]"B%�DD���hQ/���ċ��X�Q�Hl��GZ��vZ���];�.�r�Ν�����o��C;�D��䜛n%�Ԧq����rR<�pa$��AP��B�a�pH5�7j%�c���M!a��Y����Tg�^|���i_������,�6駰)�HuI�m%;��6�M�ݷ����V2lk�F#I��ݣ\�"#�#��U�`�7O�#�����ݦ���l��)˝���KOҌ=i�@��49�[ˌ%�h���9�l>�~h���3l��Ls1��y9��l[{� ���~���{1��00���cc�{�{�{�{�?c�?`� 8��8������	`��`c��X)*$s�<�s�<�)�FO"2y)fR˜�9.�.z\�������.�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��uR��K��U.�]T��uR��K��U.�]T�y��4*cB�*]T��uR��K��U.�]T��uR�B�4*cB�4*c����Ԡ *s�� �� ���y�2�
��b��cؤO�>��}}A�َn�rsA��'4ܑ'9�9͉�lNsbs��ؠ��66�l>�P��$X�
�
�
����(>�m�f6��sA��b��V˝��n�ۯ���1�~�?s�\�W9��ܘ`�����ȋS��"-NDZ���9jz������	��	Sa�M�4�(i��BPؔ6%��M�m��M�M�	�H�6�u�L��x����@?A�|�y�M[�޿-����;Ȋ��
��)��8z���AU�ay�F��NF���שiǩi�3���`�tl�W�H:�r:ȒڏM r�p[��f��[�սcxtA תQ5�
&��XtD�:"WW5�c_V5�a��6�}�ki��ک m8�mL��Q���b���mF:�O��Pq��|Y�,�/O�2��L���)�:Ʈn�������)�6����)��V��j�Kl+I�7�1��&6U�����~�&-	��a@�F9'�Ɉ���B!���""0�	�d!�m��<�q�4�r�Q��j4�#%Hաr4aH��L"F��!�<�+���e���T9�7@D��|L$�$6u���0jH�mK]My�0�P,A@�]��� ���X�Ձe~�ƀ�|����Ê��WY���[(��|/��䋬:�8�u���F��&�_��a�c5%�(ZF��`���KG��Fk���o��;/��&�DBX�f�p�LR)������q�"y1f��-�|4��~F�k�-�h�f��Q�&ԂgX�Z+R���x�ςp�rB>A�,^C)qTr�JOC�,����Y&w<[V�hYm��d��ڋ����-x�G4��kJ󘁈���S�N#SnH�sA���Y8αHֆH����KĄ�;,K���i�h��@~�Y=5�"*;)RB�D��:�@ѳ&ﲥ
{�u�����B<n���j�>��>�4���v�ڦò�ї�4�됫�f7@;
�*-i�3z�}2 ���{��${諳�����}~���c`a�1��00� / ^ �x���`� 8��8������	`���9r)+�K��<��Ȓ�*JySȌ�@�Y���&R̥�K�(�Q�ч�OL��=2zd����'�''''''')UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT���U.�]T��uR��K��U.�]T��uR��K��<ЃB�4*b��K��U.�]T��uR��K��U.�*cB�4*cB�;;}}h	P � D������J��Z=� H���������^����	�o�[}b���X��s�
lPsb��ؠ��66�l; ����(>�<<<A���l;1���Ý��i�ZnTŶ&-���i�Zn֛�1ژ�Lv�;Z�v���Ɇ�L7ra���0[@�9�	�0Na�s�`�ƪ��:n�0O��J�*lJl7N���T%M�CN&ّ7XF�n�[�jd��6�`�U�MT����6|����3��ȗ�T�[���cԢ�(�J�`�y�'��B���H��0c��?�����;��5Q�W=K_�Wtj�7Y "l\u���@��s�IH���.m�������[�H��F$�GDJ#�'Sz���A�tc��u.���k���+S��:1jעo��#Z��k�$�*&�*��J�5u6�����|j{_�/A���䙤L��V{u���f�7�Ym�bsu�\�f�'�Y��S[xS�$��59Kl�ۯZb0��%��Ibj�X���D�%��	�KBqRМTJ'��O�YМ:J&#ID�i(�:J)�
BkB��9H��P���DH�aH��P�'>	���A�&9�I�o84��5*W��M�UXj0_���kM�ڦ#
e SC�?QE�9�����zZ�+�p�ï�&�ޚ��x<N��JYR8��44(�wH�oM��
�:��-��;:�愀4����\D��M�,���T�T��J�x���A����rԤLm�d��MnHD�4�۔�jbYd$N1�&�`vZ��cU��`�{{}8\����?��(|8����8��Q>�!�� �+��p��D�B��sJ󓅃�XAV	�
aRQ0X9)?��k��;�_����>%5����X�oE���BC6��m�����u&������u�G�9���ɇQةhBL��x��
�Ĥ��V��\m�j%��
h-�����d�6���R<J�ՑmN[:�'��gu�9-d���fD��)Bt��~@��E���m6�B5��pV����������)-=���?%�2�vG��܅V�.r��cc��=�c��������"�C ���2dx,~2��, e��C�%�%���3f0̹�s��fO"2y�Ȍ�D�*	R��*R��=8zp��C40�Bd����'�OL��=2zq�q�q�q�q�q�q�q��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��UR��UJ��U*�UT���hh�4Z-��CE��y��4*cB�*]T��uR��K��U.�]T��uR�B�4*cB�4*c����և�ր@��%O��>�T�����'�� ����o�{~���}{�����; �삃�ؠ��6(9�A͍�d�(>�A���OOOl;1���ónV�������+l?NA1m��+e��v�ݩ���:c�1�|�j�ڮsw&�0�Ɇh-�`���'0�9�	�0NcUn�[��L��	SbT؛����M�CNDݎ��|�#U!�	�6�`�U���n�x�!����>A~|�~�A�o7��ǋcŲx�U�� ����$>��X<|��c�1��x�Ր�<�h*O���Ң��1�Z��՝	&�)M�.�h;7�Mm{B��\�k�-Z�ãF$�i�H��D����M1D�b����ډ���KHt�Z�E��[ۈ�q7�H���-ꥫzyjthi��Cj����@�qDm.�6�u6�M��a�b��eXw�,���B�� ����L���;�I�_Re��	���isu�ܝcW7�5��MNu�S��֛�j�x�O�Sta4�5*V�L��i4�Z5*|JҀq����D�%��	do�q��&�'��^��,��L"F��"%iHM�K0&�#
i�c��n�)�8LI��i�u�+@��&i(%M�s`�Y�Yw7�]e�RF6ϝ�>_���t��H �0���C^$�raI�`|P�J'5S�˱�ѩ8�L;4��c�\9Z�����X?��x�>���|�Q�J� ���7��L�4@�kH7�rԤLm�ĳYX�O&����I��m���Y��&���䞰S���"�0%��ƙ8�mCq��H���H��f��jJ�ݩ8HAUhI�jk1b��>%B����ZY#�PrȱhV�F��s��m
����k^/|5�S^/Zφ��S��m�1��Ѓ��%�6������Z�$��x$!y� ��^4+�B�)� �o����|Jo�Ħ�*�X��k��%�QL|cB�9�Diso/�A�p�Y>����ބہ�ts*{�KP'��5����hkO��t�9���5�F�!,V�JF��	��`��k���9=�vvN{bs��S� ���إ�C9\b �G@: ������dx!�C/���/�/� �@�c�?`���h�e�Q˱�a��1�e�K��9.y'�2y'�2y�PJ��P<y��0��<��h@�ǚ8��'�OL��=2zd����'�OL��=2zd���UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*��UJ��U*�UT��UR�CE����hh�4Z-���4 Щ�
��uR��K��U.�]T��uR��K�
�Щ�
�Щ��ʟ]�>�*}vT����p H�D��y�͡��S��'�Ƿ����������
�
�����(>�j�ڃ�A��vcaي�ڃ�<<=��r�ܭ7+em���6S���7S�~��b��V˝��l�����v��1ژ�Lv�\�W;U�n��u����nn�7N��MӦ�֪��:n�0O��J��ġ���ĩ�(nȏ������*T�j��`�U�mV���t	�H������w���>`V$oj�ڴi��a!�6Q�Q7Q�.F��F�Q��m�e�onަ�,t�),��e�%�S"Mג ����Sr޴)Z��&�RկD��5�(�ډ����{H&��j�&��}o�x����x��-�"��-�"���`��	���c�4��4�ĚAj֠�5�$���R@�y t<�kҨ�օZ��mZF����*��q|j�5#�W�������1=� �eg�	M��SvI�\ׅg5��&VO^�³e&VLp���%c�L��S-x�^b�aL�S(���Hդ�%i4��PM(FL���,��M0i�5ad��57x�L�3�����14�&�è�	xjOZ��*C!6�Mj��"�Op"�[B������ ���1�"��:�q��:�.��f�S�bM6����i|�":�L9��$�1ֵS(�
W��p��cnku�����I 4�"�ԤNZ��k �5DB!$I�ՙX��4�NœQ��6���1�YN��5�YZ� �ڲ)��D�KZR��M�^V'��fZ���H޽D�8���H�����-b�����;��
�B��F��h��օ�����!V�C�Ƽ<�k�σk�mz�u��-�x�,|7��c|x,B��$�/���S��#�S|,S����S|�<T���^Ґ���$x,^���B�y8����N�!���|�!��a�����#P?��:@t?Q#C����r޾u��&����0|�s����kĘTOy:����ܬM�@�J��V��)��8�ZVIbm�A�ab�o���j�k�k�j�j����[~T��ж�� b'�t@� ��t #�		�2�2��}G���Q���x���r�G.��\���Ke��0�a��4s�s�s�t��e�˥�K2�e,�ZT�%J�SȒ�D�ySA�M�%<�����K.�],�Yt��fOL��=2zd����'�UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT������������������hA�S1R��K��U.�]T��uR��K��Z1�S1�S�"����S벧geO����� ��ʝ��9�\�	s��'��A�����s{���=�88=���P}�>�j�ڃ���ój��x*{�=��[cem���6V��Ocu=���&( |���9땲�l��.s�9����n������kU��s�\��su����nn�7N��MӦ	���|�BTؔ4�P�`�u�m��Ϙ:�@���l�q���C����!���H}$>�I����e�i���2�?�H��C���2�n�H�ae����(7W�*$L\<�@2�7����>���,KPkH�	�'�c��8�3|d��.nSH��DJS�$�^�"ױj�֭�D��Mm�t���{i��5oV�SV�5H����oi��ok��ok��ok�`�1J�b�4ċ^�񯷇Dâ�z��M*o�M�z��: �5�F�A�\�kZMkC��2�kL�ᕇp�øeqd����4�WA/�.���%a���YrVS��&¸��_�+��u�i7p�L&�YX��i(u�Ja7�XM�V�ʞb��L��V0x�ڮ��U�V>W�)3I����p�[���=�׹�T�Ye<�5�6��|>�����Q��$�,�W��X�3�zjV�qZ���1������(4�0���G�X�x:�$#��0S�ɲ�u��`�F4O:����{nBFūr�Y�ByI`k6+�&�"o
E'4��+[��X�L%�A�t����ZBa1`S)�&����ړ�ּ�ަ�f���jkHF�h\�Y4�ga��R+ɦ"y,jhnJ�7ԫ�2�5j�D��K^֘�P�c��������Ʀ� ��8<a�xb	��B4�^u��i�|�:���$#x�B#��Y>N��M֤<[���*p���u�ňǐ��$�$���h��
+T���~/F8ĥ�Q��(:�(�p4����kk��$�|8o�C\�y4��CJ�t�� ��I���p�)b�Q΁��^9Id��w
(��A�R�$��98*�4�I�a`�d�)<��!��%8�*����D#V��F��j5�����k��m�0�!�1W!W7�f-�D��lP� G@: � ��t#�#��^�^�^�^�^�^�^�@��b9v8��e,��\0�0a�������s�t��%�K��K2�e,���@���D��$��%J����e�˥�K.�],�Y��'�OL��=2zd���UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�A�A�A�A�A�A�A�A���g��%�K<�y,�Y�4 Щ�
��uR��K��U.�]T��uR��K�
�Щ�
�Щ�^�X�����'gd@�0 `�׻����Ps}A���ou����'=�9� �P���X����4�1�	�7�M��vcaي�j��=���O}�S���u=���7Sؘ��b�	�&'�n��l�"i���vcu��	�H������Lvbc��~����nn�7N��MӦ��t�t�BZ�*lJ����(& D���"3�Dg�O��.>\H�TH�DF�#L��H����u2:ݎ�dm9N�l��q&�I�L��F�#��vD�aN�i��r6���¦������;Ϙ�j��;Z���)��'	*)	.6:juN%��: �oX�oX�MV	����[�xtb����KHt���oi�ããã���t�[ۈ�q.#��t�����:V�`�ԩ�n�[v�۷���:V	��5X7�X7�R��U�`��ۈ�H�H����E���+xtJ�5��h��ڎ�6���d�jDj �m^�CS�Hھ�N�#S�@5((��ݦ�5��V���n�5��Sqܵxj-W�Rgr��d�xw0^Z������_[���u�V>x�O�ed�q�A�mNp�[ P��z����E�)cZExm*W�-�8�RC��A��Zq�x����/��"�X׉��5 "��6��!��ʗ6���o��!�������]KV�"�o.��Li-��"o�usn۸Vk4��L�Y��n�E��n*�h�����sΐH�Ċ�ĥx,�k�1�X))M ժ̮�q7+Ƒ�I��5�E�W)T��A�)����C��x�v�y|�j%�Eh�u�M�>=���S%��,�'����RQ&��<�R\+�LF�w���M����Ag�&�p=@U������� o��F� �	�� �1�/x��@���<B��(�_���B��SI��ť|:�����?�����B�y�����j��JJIY�X�w�ۃ|V���:���"����~�w<�$��V|�Q%��ʑ�_���9ܦ=%T��mz�#�r���p:!8HDbN�#VY �-<F�#P��O��*��m������L}��L}��L}Ƿ�=�0: � ��t��?#�~GD b ��c�8��Q<��ȆT0⡉Q8�IX��,[������9�9�:Z:Ys��%�˥�K.�],�ɓ��e�˥�K.�],�Yt��e�˥�K.�],�Yt���UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�US�g��%�K<�y,�Y��g��%�K<�y,�Y��hA�S1R��K��U.�]T��uR��K��Z1�S1�S=�������� @�5������	�o�9���	�ou���'=�<	��P��$�S�S�S�[v�ݰ
�l;1���j��Aڞ�O}���)��{��n��1A�?l"LNT�[\�rD�sA�����4�7_m��u�����f&;0���9������t�t�:n�7N�6%M�CM�6	�P"n�"L@�1qb�4��M�DM�DM�DM�Dm�Di�7XD�au�m�NDؑ6$M�CbP؎�#�8�N6Ӑ6d���e�M�6Pi���lI֜��"L���Z�ޚ�����$�h'������*��㢤�����.&��YT�J�eH��#^��ڹ�MR)�H�֭�: ��5�-Z�-{-{-{-{-{-{-{-{GK��q+��MT��n�[t�`���`��[�emԖ�Imԕ+}R����M\I�-ꤊi�"ޞX7�����E�.�k�֧AM�^��5��h&�}i���m�mS�F�= jPH��Z��5��#Z|�kO�F֪���QZ�#kU�ڛ���U��Dڦ:���Sj�u6��Q�A�:;:��7S^�k\�f�����a��5���=ӽ2{�DE��Mt�YL9I��~��������#n �@��n�ʹD��Ÿ7�H�$F@���_#s}\-�m钔bR�pn/:b�y�%��f�W-rP�u�Õh��p��S�qy�qiZ�:Պ��x�>�����:ժ����jk��D���W����m�&��|v'��SZ�X�_4��r��H�U�W�� �R�^!qr@nn��
�'����c�=DVmI�L�m"0 �,B����B���b��zn�a��oC�d^,Bk�7�x@�Bi1�����?�7[�,�w�׀aU��<�w�_�Q���x���PbLl��W���B�w�����q��W[����o���u�C���$Ғ�.�R��JR;�JG�b�������\:�(頫�y��f��H>���~҄W����53�"m+[��X�	MBu�H���$w�[����:�N��4�[�GQ=0@8��f'6�:�5�n�tj@yH՝ǋ��<��#Z�0P�>�ߠ�ӃTTS����'����T �t #������:'�t@��3 e���bTE� d�!�O8�a�������	o�(�h�h�(�(�h�h�b�E�9r(�Q��1�c�`Ìq�0a�8��],�Yt��e�˥�K.��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ�y,�Y��g��%�K<�y,�Y��g��%�K<�y��4*cB�*]T��uR��K��U.�]T��uR�B�4*cB�4*``��� @ �{{���^��A � � � � � � ��Al`[ ��
�
p
p
p
p
s�9��{��0Li�ce�M�ÝAڠ�l9�nV����n������{��n������{�l;1���ó�l;1���˳ �7�M��}�;11ى��?s�V�j�1��ƪs��j�1��j�ک�u	�b`Ӗ�XT�@���Bb#u	���BZ�*l0��¦�
h	�(lJ�&	��t�>T�-P�-���Q6#��5�*N��ʓ�I�6���!��vHْ6bG�m��G�)/��H��D�$F�"
e:&�H�j�.H&��ʰIR-�j�V��j�\M�"��SU�j�o�&����z�*ʥo��!�RխA"֠�: �oX�: �k�7�j�کjעq7�R��5�f���E�cxmc����U�Z�֤�Ԗ�JWy\GDF�$֤��U*j�oPH��D�S��Z�R�dХo�8����"ޣ��B�M��~R�����|	J�}q֭jsxֶ�b�Qd��mLá�ս?o����Dm0o���e��6�Fè��u6����NZ��:���Z4:�����n$!n)��>;#���6��9,iAr��&��9ݬQ����/!����x:ۃ�-H�jb��|����ہ��'�[��=�4-�
b;C�V���M��G.�[��r ����BS4��L�Z�Ɏ#�5���p�xM&�%"��`�x$����H�N$cx�>�Ui���4�B"�D�V;5�yH�V;�f�aX�M,�
��ݽ%���խo������w!'��s8ǋnRZ-B�37�[W��y�`D�>nX^������Cn0�~Q�w���!����D���������	�ǂk�&ҐF������H<�_��Q0��l:� �i1��H� a�[�^�z�_���������������|�_�^�����A�c�^�pA�Bt��Z��\k�|�y��&���i_��h�k�K���<���$�\CMo&�b>Z7��ٴ��)7J�y�s�(�^c�4/�d�ʜX�y�v��PN���@�19�M������׉�q��j�{M4�J����|��*n�"O���
�69�'*~Ks~�3G=[}8	�p'������/�]���y��G�"yp�ˋ�"J��	uQIX(bN�31���oǆ`ƈ����
3��r e�a�t��e�̞�=2zq�d��XÌG2�9�at�'��O.�]J��U*�ƆhbUT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�A�A�A�A�A�A�A�A�S��)NR��9Jr��)��4 Щ�
��uR��K��U.�*a��Dy��4*cB�4*cB�4*``����@ �{{���^��A � � � � � � ��Al`[ ��
�
p
p
p
p
s�9��{��0Li�ce�M�ÝAڠ�l9�nV����n������{��n������{j�ڃ�A���i��o��+M��}��i��Lvbc���j���NcU9�T�5S��NcU9�T�U>�O�S�퉃NZ�ake��4��j�0�m���Z��R�"�EI�'ʓ�I�(0M��CM���S幂|�>:�a�A���['�4�9K\�mڜ�ޑMH�LzRw��	�b��H�[}R���v���M*5��,Ԍq7�񽴇Kn���*�Oq)+�J�V	���b�cmԖ�Imԕ*ʰMR'DƵq�O6)�e=�X�jJ���Wz�+}R�Ճ{q)����5���6�,�T����e5�m�Z�L����	�%6$�e=L���U3�ltV��*i*�4e�ޗq&�8�C!K���^�kݒ-����kܛ�jsHڧ���5���ֲOY��$�ejtLo���?i��*�=�mn��F���u�o\�K'����,�5%bI6uU�\5���WG�[�:�/I���3h;���&6�SP���V�
K(� ����!���ס{���[�:�0�M�Bk�@�H��d�I��H	�2��D��GL#Ջ3b{����4֑Y����$RoAt������j;��Gc��j�V�V ��E�k5�T�W�nۿ͆��\��+��A jԤLmͧBa��"���\�i4&�L�B&��D���Y9����;�� kdU�:����!�t��$�ۈ� M���jm�\�Ł���:�ͺ0�׷�N��Jq��MmP��T44�o��l:�m+R1��7-H����u\H�+������ �$ǂ�1 �LHX�8@�.�����i]n����i]n���/x��������c��/t��Dc�(�t��@u���k��&�Z�q�N2SեZ��1��~�(�F����%`�rﵦY��xNo�I&T�I!c�Ҿ�g�� :�@�� Z,V�nx��-1�J3�N��)%i\�"b}S5�#s�p��������Ƽ�Nto�i�۶�����DbX�#O�Ki�bp"��7b���(A�,��$t�J� \�8�ЄQƀ�җ<���T�Ъ\���-�&Z�e ��G9.z�f�f0�a�t��e�̞�=2zq�d��XÌG2�9�at�'��O.�]J��T�C40�C��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UZZZZZZZZNa�,8e���2ÆXp�4 y��LhT�K��U.�]\��u�S4 ��#�hA�S1�S1�S� ` �} ���1�3�1�3�1�3�1�3�1�3�1�3�1�3�\�V�V�S�S�S�S�TX��ƛ�74�P}�>��i�ZnV��+ll������u��l�[)���s�<<<<<<�
�}��m7�eٍ�f&;0����U��h5V�j���NcU9�T��O������U>�O��M�'�s�9�#�&91�����h�0�9�I�	�."l*"l*P\P�\n�x�A)�z&�s�W+U��}�Zm���5�I�7(�t��I5jf�s��bկD�5��F��#j��ډjmDhII�(I��5Ј��DOS�WX�jJ�eoT���RV
Kn���J�Hū^y`�\kR[��ֱ��6�O6$���Z�x֮i��F���kZF���k�$[�4�z'Sj�|YJ�4�WU+T��t�SV�ک�S۔��k�)VWi���^��6�o��S��z�`�\�X��X��X��X�m�-���n�<kIn\K %��H�R R��M�$����tsR���M�կi��ke�k�n$�{n�rY��TMkM�֧�VO�ˠ�r�8�k_N��R^,]!�D-��Ӎq�8�^`*Ȱy������~16Õ�l5<��$�1��M\S!��MH"�t�A�!w5��؄,!|����H��2���vh^�AW������ʈm��:c?���Z�+�����$�M�u�wZ��$��� �%, h5jO'���PE�n/[Sx?ۋx�>	R�j�Y��k6���R����`�'��'b{H۝��Sb�ĦV8��ũ�|�m�cSI\�S'��sU�D��LBn�"OU�Mppp��o�[�h���� ����8�>m
;�y�j��v����pN!&���A󈡩$H�&�����Ad��F��$h�HuU�a5qм z� ���1x<p��$ę ��</p��#��[��x�ŏ�{��w��+�{��/x=B��Q��
< ��Ǩ�I�w���6�Z�+D�d���$x�8�k'q)H�>��q"���[�Ԍ~^7ݦx�c�W��"�<
�P0��#u���Pc��FV�!`�bp���3��j�ܡ�5rFS�K�H�7Z�.�u�т$ę-��+(�@M�#�Lj?Q�GrZ�<un�#E$��ڮ�!���#��*����U��c�E�c��q�]*!E�
.�0dɘ�� �P�ʐ�"�GJ0⡇#�\0��3^\�a�t��e�̞�=2zq�d��XÌq�0a�K2zyt��UT��UN40�C41*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U�����������������2ÆXp�a�,8e���B�hTƅLT��uR��Ȫ�Z0�B	O"<Ё�1�S1�S1����4f�A�3_�����������}~��]�1�3�1�3�1�3�\�V�V�S�S�S�S�TX��ƛ��f(>�j��aٍ7+M��r�ܭ7+M��[���7*s�9��
�
�
�
�
�
�i��o�����˳�~��#�&90�ɇ�L>ra���t�9���n~�?[���ܩ���f&;11ه�s�9��ܘn���
�	�.P\P���m��u��u��s
�����̡�&� i�F�r��O+mɩ�O:=���_u5�S_Q7��������vIVJ��@ز<۵�C�@��mQ�k$M�B�ڹXtD�&��YVkr����q�ުm�ꕾ���7�F$SVݾ�Z�8��8��,V�I5���J�p[u=`����H��C��okT�"�V�}�k������WQ��hQU)T����o�&��YT�n��)*�cnT�Z���:%��Sn�<�S�m�#u���N)f�GnT�浈���J�?)[��;�H��;7�{�Hק$��&�m ׹$N�T�:��J�8SOW�Q!xD���ǘ�+:F1�@��Τo�U��:��Lu7�3�ވ^%ԱW�������_�����i|�Q�^iZ��Ԟ+UbiD��|�{W�c�u�ŏMZSp-��d�p�^``��)�f�h�/�ZM�8�w��A|�'$�e���׵�&��'M�"1�")$I�5�,jۓ��RY-�4�M�{^":&�F�hH�w	�@Ւ��ެ���h�ڦ�Ƥ�5�o����4�t'LD�x�f2r�dҸ�����=U�kA�T��������Đ���-E�r���pc��~Ԃ�F��'R@�_��C���ԚGx��>u(���(	�����۵[KxD47�J3HF�4�`D����+�eb4 �/����4�ď���/��L�<�
��Ŏ���@,u��������6!�G� Q�@>F���s�y�F5�1'q(&�.�
1��Z:�:��n[
#����	�T��t���C�L(9/�ŏ�0����p�������_	��B7�5�p��E7X؅Z�Q�H�q`P�<X~�-�E�M"T���7�ɸ�H�bup�8qW)�"MDML�ߞ��QHM� <�#hI�r9?_�47���������@��4.�]{�d����������� �� ҀGJ�qqt��ˢ��av/20̺Yt��fOL��=8�2zd��XÌq��̞�=J��U*�US�8��'�2y��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UV�փփփփփփփӆXp�a�,8e���8��B�hTƅLT��uR��Ȫ�Z0�B	O"<Ё�1�S1�S0 �P�o�{~c��@dE1�SE1�S�1�S�1�S�� A�3�1�3�1�3��ou���'=�=���l; �vAA�����ó�l;1���óvÝ��l9�t��p*p*p*x*x*x*x*x*��`�������/�7\�?s@���4��?s@��~�?s�;S����:c���n�[�����n������kU��r���Z��jz	�0[��O�����*P�'D�"M9#��Ӻt�vb$.�)��N�F���"Sz�ׄ��������;=�d�P4PD�]hR.����s�w#b�*@���,��w� ޠ�:1D�cx�\K+n���5��kXە<֧��*ս�TƤ�tN#�`��u�f���6�IH��$VH�������T�k�u*ƶ�mk�U\w��H(�ڹ�T�6�iLH7�4��M[���MV��վ�VV�cx�1�Y[u��R[u#�DN$�U�hcx�~H���!JU";n�.�YR��8�CI���:�b]�I5���n��WH�H�8�6�n&�АZ�������Ym�A�6󬗯:��Q��L�ͯI����i�^/���x*�%�J�k�9H�G�z���P�4��P�C�m!���X$H�ܚj�2�D5^�
�#���惡!C�C�/��@��Gv�L'�6˴?�K0���N)��&��^ވ��hH�NR���h5jv+���t���+��D�b��LXF��Q��j6��%��L�v4����H�V;����1JW!)N�%�rZ�� 4jWX)�@A����Y0�V4�=sE:�@�Ю�ۃx�Jā�bޒ	��%���ư9Q�H0��r����6��
:�������ۉ�!��ܘ���5���Hѡ``.$KZ�����J�e�@�*4�O�@��u=�7��&�+
�
� ���F���©20�L��I��Rda��y�:,u�E����!u���У�>x��$�� ��H�k	N�bLl�8I/�����h��Z��Hk!xH�#	��a�r 묈F�$
�����0cĠF��G���W����F�JƨU�Fx��\$AD`���/���h�|&#I��у�X�u&�iB+��o���	����Ҏlj�N��2SZ��N��\B0Xۣ���fʸ.Pi�i�"�K!�����sG�3r ̈�QCe���^�*,�dv�꧗K�`�tINZҙ�3.�],�Y��'�ON4N4L��K.�],�Y�Ӎ��UN40�C40���@����UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UZ-��CE����hh�4R�A*T�A*T�A*T�A*T4 y��LhT�K��U.�]\��u�S4 ��#�hA�S1�S1�S#�
� *��Ƿ�=�0dE1�SE1�S�1�S�1�Sߘ��Ƿ�������}~��\��ou���'=�=���l; ����T�T�T�U�aٍ�f6��vcaٍ�;a��s���
�
�
�
�
�
�
�
�
��Ƙ&4�1���e����dI��Lvbc������f&;11ژ�Lv�;[��뵲�l��/����n������;U��r�("-P��ګv����j��V㭈��� .��dokJ�w��k�b��sZȇ��(�
��������Y����+N?��H�Y:f��7���jg��$� �mMf��,�����(.�'^�����f�N��ԕ�Y.�4���!�%0$��izł�۩��S�JJ��R��5%f���$��&'��0j�i�mO+�A5H.���mk�U�t��(9L�0�qJ�RV�eF�<M-	3R
涬:U�Dfև	�+�����ֱ��3�ܸ&����Nyf�hY���F�B�c�q���L�\�X�R����7����$)%Υ�U���Wj�Ρ's�׷���ۉݬQ�M`H�(���~�%=\o����^/���\_5�20Dn	�u=!`M�;�m��=&�t�4�^�'��^$]D���"O}?��d\�ځ�j#|���\?(�%g�TT6�S�w����7�!�,0ǽ��M+��M����&\D���6��d�ܖKm�&��L�v1I���.BZ���H�m�M�ӡЄ׷�&խ���^t&J�ba5���pi9�	�`�[r'��#Z��kH6���zR4�w5N"�E�Ij3���$��a\:�R�SC�Be�ñ�p��0�\�͡�:�`���w����l�
�3������@�;�� �pvL1��Ãn��gÃn�v���>m.&�RH���u"�4��d��Y nu�TF5a�MX`V��B5qP1|P_W�aU��Ux&^	�dB�	��Fp��]c��X���E����h��Ą(�xy֍���kA!c�V�ń� y�x��`�M�Fp��7��MxZ�/
��c��*�"	���8��DH6B��{�!x����r�H �-
��Ѱc�� �z�c��0*�+����1��&8$
��GCRu�Ev���:�BNrspY����iD<.$�	�1�Np"k%,�%���S���p�8����NLM(�M������c�<e=���ʑ�O!f)�����e�˥�K2zd���ƉƉƉ���e�̞�h�h�U8�Í8��'�2y'�.�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�CE����hh�4Z-����<y��0��<�ǘx�a�4 Щ�
��uR��K��U.�*a��Dy��4*cB�4*cB�4*`a�1�� ��t�"}��R H�G@: ��v���� 	��~c��ߘ��{~��^߮ow7������	�@��	�H6Q(A=��)�t�U�6�P}b��j�ڃ�A���O}b{��X����(>�A���OP}cL`��}A���e��&����/�6_Pl���vceٍ�f7\�n���s�\�7ka��}��]��jc�1Θ�?[�����M�'Ϝ��s�)j�u1pU�mBtbh�ڑ�-��	�+�5%�5�C����<.�I�Q��1�< n���t�:�ӏ��r?���޿�Žt�|����鳩H#�^��x��!�]�7@�h��w��>u�S�o��xD���'��M!�Wi�ƴƦ�LQ��J�q��� q�"QH�9I��MGuҴ��J��+�� �BN:��1ؔN{V�_�&��R��k��p��6�84�ͥ�PJ&�npC�����M���[Q��ρ��a��Ҕ�59' V���+�BA�D�o��Y �R"R�U)T��u�B�N�֧DkS�5�سX�۬Pi���+Ĳ(�Lr:�������u	׏T��y��Z隙��Q����x�� m@н|�Re F��\H���&�[��0�F��_����W�F��6��|J�I�5���T����;�D/nƱ����ø��R+�cHSw�2�yrԞl	��j��m֫nm��<��Y���"�D�Vm�cU����S)�� �@.H�΢xI��r��vW6��"�X,��Y�͇gP\D����!��Z��Iy1f%� �[rO%��&� �Q<R�u3n�kN�L�h����Jq=	2`ym���D��n�"Y;ěscr-��m�t�"���z�3��M�`�"��o:մML�H.$D�J���͖�Bv�m����m�q�n��thR�6���iq7_&���o�&��,�?|��gQ�Y�|u�q�A\`W��B5qP�\T_W�AU�UxDI���27��:I��c��Qh�Z^�����0x�0?��j�q�8�1�Hp��b��P��Px#_%��1�FW��E�B��F�#/�Bj� |#u��^aW�@ux�m*&�u|`��$A� u�nV?��0���&�0<Q�2S� �*Q����9 A&&�$������hi��2@��F�/� 0��� �$��^����S5_ţj���v���$[��"s������j�`V>1	
r����r����e�Ǯ@-�(�p�.f],�Yt�'�OL��h�U8�2z],�Y�Ӎ��q��d�O d�Ң.�UT��UR��UJ��U*�UT��UR��UJ��U*�UT��UR��UJ��U*�B�4*cB�4*cB�4*cB�4*b��K��U.�]T��uR��4 Щ�
��uR��K��U.�*a��Dy��4*cB�4*cB�4*`a�1�� ��t�"}��R H�G@: ��v��=�b ��o�{~��1����{~��^߮ow7������	�@��	�H6Q(A=��)�t�U�6�P}b��j�ڃ�A�����J�����6_Pl���vceٍ�V���i���l; ��M���`��Ƙ&4�1�	���u�|����:c���l>� �7�u���Lv�;Oܧ�S�)�ܵB`�7r�9H�/S��M�mS���5�7YA������S� �w�Tv�z��E��A\@I�5��1��?;�1�<���@�b��,C�Ә�w��V.��X��Z��Z���5��X56�9��z6��U��֫�~VW����=3��;��c�QG;��3Px�׽�@�GR5�Ž^��@���/Z/[C��zgA �օ�|#w����Ь|�#���>���+z�Q��d>!����{��F�K����j�
g6�~����pw,f�"iV�&�����
CNԉ��_��cH,V�c�7X�U/Z<��1���T8��]=hBsx�\�f�'	�=&YN^ܗ����R��e�i2�1FK���T`�h�T�pE�w[���d�����Iz�w���N�h����>�/h1&&u�EŨ��������_�[`������\>|�u^��ɰci�pF8���nY�G��Ϣ�m�܀B��@��$u��j90B�5�g@a$�))�WK�"�4�ڍN�#b��_-��3Ƴ�x�H>m˄�W_6�7��\����:�D�_/�+E���x�V��h	(�	RM&�/��u����o��a��R),��U1�k'��F���LOogf�S$-˨�R�T����8��H+�E����]��+�J"siiM+�.Ҽ�4�Z:�*��� 4�n'Q�ҋچ�|��b�B�;�o�mo�Ѧ_5�B�h�HW�$��*|�@���ۖ�|ܶ[Lp5��śdhmۭIJ�Ԗ�j~�7��3H�$ ��"A1�H>J#���`�:��Q�MX`�+�^�qhA|T_� ��@Ux&I��W�AT�Ux�/�T�l$#Q�d�r�H^�(w�_ę�Ux&�7��q��F/��%A�b5�u�=7�|&�8GC�����
��Dn'�xP�/���kJ9
�H�%cT:�0��ê�Ы�tX�F�Ն F���<Hêƨ���	����q����o�����"a5�S�S-��E�5�Sо0��5�h��:�$�¯CRV$��3���j����c#��]@Q/�v�y�o�Q�w�e�k6��ߚ�ȓ�Z�D����4���˜���92�d��C��U8�2��'�2yƄ.a���h@��<�t��c0��%Uhh�*cB�4*bUT��UR��*bULhh�Uhh�Uhh�Uhh�UJ��U*�UT���S1�S1r�.T���˫�W.�]\��r\�y��4*cB�*D�%�*]T��uR�CD��%<��B�.h\�r�K�1r�.T�C(c`��1��02<2< �P�_E1���)���T����������s{�����ow7��������'�A<	��P}D�삃�
�(; �삃�
lPsb���P{T����Su��L?>}��O���;MΠ�Os��_\�n�N{b{� [ln�bc��h��?}�\��L>v�@T[!��v��Wd�ȏݑ9"?[\`�������u�t���I~��4���)S��yIM�P��iHo&�"$�!�5�4k\�k��I�R�B�
:���6��w�W��6�Gm�@�����9#� ^w��n���MCppABQ#P� ���X7C�c$�c�b�7��1�י�<�8~׺`���M��i�\V&����Go�M$��t����n?5��?5�8R������?���~:#�^�-{��z�ͪ��[�Zm[�Zm[�ZmF��wB��iGw��/�-C��Lv��Lsh����?[�1!��4��K�E1���o�_��ҿ1=!h�����]W�w�-F�p&=&�mo�M�o�9��R6�y�Oy�d�qDb|�"�\W=Bo!c��B:ң	o�F���N�q_�͡����:I����GxQ&:�x&�i���!��]F��0Zq�P0�p;<�f���У5���/[`�P iKn��]k�囉�_�Z�B���~]q䬵A4[���y��ԙ�F�1����ڵ�Rk��%���tPI' \�R_,��I�J���W���j�q�IJl5��ʸ�vQ��#a�|vnU����w�-��DBX�%r�X�K&�#Q�زY��E"Y-LB!ƣSCjm&��D�q,�i1�)&�jS6�J]p�B�M#x�S�g�g���.8H@����Q&�n���$���f���B,�^.��P�W���_��(���iA���7毭�*�կ���5*1���9�l4zgg6��?��6�L ?�]�K����:�A_����<>X6�+L\mۣCn�m.&�iq7[JE1�-OƆ������K���+�5q�A|�/���T*�-���j���<�($��2��L��p�����c��<�("o�M�u�?�����T�:ʂ�����&�$	�I�0�ĩ�x�B���AxnW���A��о#�������&�7��B���W�
�ס\Z�+�^�qkЮ-zš�PA|T_���PAxZ_�ůB���V����Eq�Y\n_=
��Xn46���xF�R53�<IR�>w-���cc��;	7�\���5��32��aI4�#n�r?vD�n�O�Dғ��gB�`*�@�=J�}{2q*�L�e*�K�8d�9�����茊~���),�($ys�ǙCe����R�8�a�4"�EG1�r+"�%<q�K�y-E(!A��8��U�O"8�ƅLD��V*���Z��J��'�1)�J�*T�ǘq���W �B�� �uRY���k�W.�T��BUK�*T��r&�Ț
�C(c`��1������@
�}~��__������������.�.�.ow7�������s{������lN{bs�� �	�H(; ��{��X�����'�Sݩ����(=�P{\�{\�{A�	����i����i����շk��m����P��
xk`5��n��O���h���7A1��l��Ps3l
�]�'*l%-O@��|
T�X�M��YIm���ƅaC�6�y���h���<�%��%I�k��Z�|	���������F>������"6�%8�DMc�H�Q�a5��@9t�#Ł~��I��<���c���n"E�Sz�͡� :�O2��zGSȰ:��Ө�m
q�zm#�����M��^f��[���N�@�jm�jkLu�����t�M$�����7;�1�A���C����z8����+���o�Žo�Žo���C�Z4��h���鸵���kF��֋s�ߦ9�i�qn?E��Yo����G�˧�WL]0pmo��^�{Z��M.��6�I���I��&�S���d���zk�p�%���lc,[���o��������	�P������>|>N���l�eB�m�D�F�e���1�Km�L�-��hHg�J.Sa�߮��.������Ʊ�I��JX:�j#k���Y#Mʓ��e�*d����nT�c�/��eƭm]�ִ(�:х5�4(�Q2��˭Zu+[��u~�xuA�ge����nN�'���I�J���դZ�p��56��(�&�<�MS-R
�[r�+���iI"8� թ��'��F�jD�S;HJQI�1�E��0�K4	�s�܄ڶ� h5je��Z���2�̢����,x�Bm��+(�Ce��J���C�f�i9����B4�2m�^�~W�u�8�"�`����X�L�44qn
V��i7��c����BNkCIìD&�-Mہ4b�5��5�x�ۨM���m��Ͳ.,�#Cn�jK�RX4ړ��4$S���\H5[K���]G�e��M|~#W������T�0���j�b��0$��Ы��*�-eO㬨*�-
�KB�Ы��*�-
�KB�ЂLM�_�c�Yk��j��-�c�0 �j�K����|�C���AXF#W�B��W=��\Z�+�^�qkЮ-zůB���W�
�ס\Z�+�^�qkЮ-zůB�� �-:��SU�u���uX�|���5r`AX~Q�U�Ђ�_����Edq�j~������p�?��8Q�6��G�V��W��Zt�U�@�Il��S 8J+���6�jtcE��i�C�9T������,�&U q�)ĦC2e�R�*JйM��SL��ː��X����ƃ�ZB�1���̞T�r*R�A)�S��GDd�arꋗT��$L��Ɔha�*b�Ij���9J�y��zЩ��T��C�O.�A� � ��1V��E�J�
���T\��
� ��C(c`��1��02<2=�d2<2<2<�!PB��A
�}~��__��������09�A�`s ��� ��'=�N{D����H'�A<	��O�{��X�����'��=ڜ�Nv����i���େ�a��{�@1���l�ce����ݦ�l ���V��=��{�_Pn�"P��
���6\�&9�n����>s��H��	��� Vu�Bǫ\9w��D5h���T�?�����0ݥ|���T|�-�B�YP��T�Z�G$N5���h`�!�4��6��T�V��U�B�u�Z;��C�h�U�&!V���:5�������%x@w�O;������hw�����ā�F)�ءhRn��n�pE� QąӨy�@oIGy�;��Qǚ���:���p_�����C��1���q_�c��鎷��:�H�p=&�zM�N�ε#�:ԁ�֚N��ru���d��'�?���c��H:#�W�;^�3��ji�u������:M�d n+!qY6�M4�6�ȁ�]#��際ZX6����Z��G++�zM���<��P���3նjoW�$Z<�o�����-�灀Q�n0+KG�����d*�n�u+�q'�N!ШD "�8��X?��[^�J4� �F,w�H]W���V���m�bH$א#\�73�g��J�Ѓ*Q͊t�D��$͡�j�+Z�;z�/�i5 o\�� �<@��I�S7��1u)d�N&�Mzh��I�f�1d�W4���sB��Z��u�	5�x4.BZ�K'bY��N17$³rR)���)\D�7$�R̮�owZD֓	��ɠ�i;
gbid�S4��D��$�-T���~<�0`�xW+6����xڒ�Nu�Rr젉�S�%���5X�������;ί�c��|��У:McP��Ӧڂ�9/F�o�ӿ��ÓZ0�:C7y�h'�r���y��Q��*p��szjd��lP�ͅ~kl>sZx�Ot椥O
I`�jI�еn��"cii�e�YԘu&��b`MX~�+ޅa�Ь7/���TF�7���3 bL��0$��3 bL��0$��3 bL��0z�CH&.(���L��u�g�4�T,�*���>I���� �-+���T&�>z�B���_=��|`�/���о0���cT:�j�U�P걪V5C�ƨMDn�4��CHZi
���Ң7:�������/I�F�xZ47�A�DL~R��	 �X& ���_	$J�H��k#�^�sU�ޣE��k�
DڶMM�T���F�kǞ�S���*�S���r9����UTcD�+��ȁ9�["[����l?s�
�9Gh�K?rTP��ȼ�̊.�0��Z'�E�9i���=�2f����+�bSȕb��ǘ��J��U1*�\���%Dd�	UW.�]\�8q�Ӎ�����A�"�V��Ɗ$��g]s��T��.T��C(c`��1��02<2=�e�d2<2=�T�!PB��__�����f;c�f9�A�`s ��� �09b�� ��I�lN{bs��؜���'����>ӝ��t�js����
�	�@����4� ��c�	������ 纀`1ه�H�ӕ'�6A[�h�*n��i�.O�x%����5T6AZa�nU�T��T�6�jjV���*
�	c���Ѝ�x�B��ȱX�p��\'�G�dB�i�խ1
��B�7�
�j����X�7+J����\~�V�&ֆ����J`�#����8��>x���4�P��P�Z$O3�& !���� �]QǛ����ƅ�#�i�r����-k�u"�" y��'�m�y��b��Cѭ@�t@�5 Q�
< n�1�$�6�7I��M����V��偌�,C��m�t�I�2H]1�N����3qt:f��t�M$�ښH9jk婬C���t�R��:��ԧy�B�@u$�RI�:�M`N�<�klk�����w+D�e��@�y/]`n����F���)(�BJ0<��1����"
��%��ТO?ς	6贳)*|Z���P���2�^��8�k��Iz�o�٨ȷt��@���7�<�CpZ(�bX]d@$�7* i����l!X�����E8ف�O"A����4<���L �oE�ƽܭ:5���\m%���]u*�H�Nn#��F�D5kIm����:�����2�����;����&�n"�h�q+]i6���w�Sq,���S���Pq�Z�:�- �&��.��|�w���!�թ5����D���"kI������`�q�H�m��3��ƭx�Y�!�`��%aM~]�'7S�/:A�,�Z��B�iܖc#"���5�&�`�Zo�l�<���_8|,Q��̣N�?�-�0X�R��^�_��Cr�:�nF1�����!Ğ�?�B��vNW�e��kr|�7a�J�4)\ڒ�lhq'	�RZ��Kx�Q�F� �|�����Q6B�&�uԘu&]I�5a�Ю>z��B�� �j��P���_5B�A|�/���T �j��P���W�w�~�-Q���r`1&����i3p��?q���-4��C���W=�M\|W����5q�M\nW����5q�M\nu�G�gQ�Y�|u�G�gQ�u �	��5�k�����kRid��MD�(�"���uj��5�0|��`D���&�?�ƅ�\D�$
 �"7��	hM{��`HBtp&VMY����F6�1�JY�M�:edoXۦ�SMdT��U���4�6ؑ�I�6E*���S�]�H�憴��ti��f���v�1�}i�����H��#�Wrb=ؼ1�U@Q��x+�kM� ���aف�L��ET�*�+�%AZ���ӈ��_�C4QЊT�IQ<��TK��'��%�=J�yuRȨ"�VѪ�+�Nat��Xʦ�LA���+�"�0P�
�C(c`dxdxdxdxdxdx!PB��__��A
��__���`�v�`�v�`�v�`�v�`�v�`�r~A��'��1l`[ �s�%�-���������������\�\�\�\��ow7��� ��da�LL>~�CT�'�\�����6�7����h�Ϝ��[\|䉺�l��;0�ɍ��ؚu�a'8/��c�xZx#B���bM�/p�G��Q&�Ҥ�n�����
/"��`^�O<������<�ǉSRH��Շ��[TX�>�!G�a�F4��v�\�>i^�s��6�>M��;��A�Y�xP�/��0��|�����~�>څ�ky�PqЫ�~8(�$���ۛ���W�y����4kP9k#��QlJ#j	DmA(�@CF��4kP$jth�
H�(�n�p t��:���po��I�� 2��z��~X7��u<�&��6�7I��GS԰:���p_��;�]���*���W���]����W�`E~��K���@Jy6ġ�r�u�Z
;����o��|�(��*Ѻ��(���|/p�׍���@�l�F��ܹ���֦�L�A&�������w���������\!t�m�`�7��(��f9���d�a=�;��F���4:TH���E"/4�n-�,u$	����'� � �rO-OBMN/F7�7��|�R5��K��)�֠ӌ�8��V)�Z��sU���L��nqr:1�9W�R硩Q�q7�4#��u���)Zu��2�u���V���;��%�O	&�Z# P���n1�1���|�Ÿ�q��5'�#zf;in1�"�1�M#������\�*>j��n���$Ӹp�Y�
�{RH��i��Std�C�U�f� u7"��5w�=O��\[�~7�,`���m-�|��b�~4>A�~�_�|o�c~G�.�p���U��&�� �WN�t������� ���'`���-��;r	�/b�� �ۀjJPCB���,��sRH�������6f�i`F��H6%M�Q4�%L,�l��M�걺V7Bj����0&�L	�����о?z��B���_����|~VM��0jKS�0F�n������*�Gϝ"�m-�Y nu5^�q�M\|W�MP���u5Bn��M��	���7ST&�j���d��Y ~H���d��Y ~i�m�T&�>M�j���&��FH�M����u4�#a�ogQ�Y\n�]Gϒ�0&�j��"c�*zBa�	 Y�*+�䥊�H�	���j �@�4��19���xM�6���!��d0�S8J�eb9�N�0�GP^�f���i̲�&�n����7�k����xjNp�Zi��x5N1��R�|�Uw�&�F�qt�V5����#����fF�ht	�&"_�k@��$f^E	G��uPG ߏZUDĬ<�2� �8�0T�����K��NR��=hh�98���yU�r�%��ʪ����ZF4@
h\Ѵ1�C(c`��1��02<2< �P�__���`�v�B��__�����f;c�f;c�f;c�f;c�f;c�f9�c��9�c��A���`[ ��f9c�k�k�k�k�k�k������[[[[NO{ca퍐l�cd$�L ��6\�4ݒ�>�NOPl��CO�O�O������P�8�b&�pI�s��hq5EęPA�`,>
�����
��|�v
/�T��J�P8Zc��x�,p���`��pA��8O�i3qi�vQ�F�1�|p�C�4��=�x���i�G�L(�i���ź�F��Q��,�>	�����U��&�6���^��`u�1z�*	�ڒ@�qR�-J
��(q��B���l�j�i�q6���V���2�M�|/_i�P�l�&�!�5�6��"m�r&��"j �mC΍I8؁�y���0y��6�Q��
6�F�ǜ����$�� �r@�G�b��r@ %5�B�h@�-��l�$t�H֠�F�|&քmaI6��F�/G�&nu�ъ�t�{�8<�l�͐��@?R��g`M�L�1�e������`�⯃�~�E������y�e�4���]0PX!��PE�:�m�A~�X�	�7����M��`��[t�Tri[�n#M��d���4� J����M&��V-+�d/x,B�P~�mZ��f1��D����q]�7�����n\M�� h;,m���vo)�nۯM�M�Z��ł�LhH��F�x��wkI�"qخm�D㰈�v5��ƑēQ-]n���D�u��W
MԴ!�[��?�o;H�u�����S�$�L���C��sa�m`!]F���;��!�L�5=F2y���
d�MhS>
aݯ1	6SC��&�d�_���"�|�c2	�^� T ����8m"�� A��6��Ö�6�B*ӳ��<�5� SC�������a��?�=2{ڿ6 |��Á��pY�wᡷ Ԕ���+�RX96�sRH��$�{iZ�6�����((�"r��'(�"p �|�M7�D�|�M0���u6BΦ�Y�����ct:�n�U��걺V7C���Y�|-,گMJnԖ�W�D~V&�Ɂeq�XZ��-P�jn44��ET&�?	�����YX����#���:�>����#���:�>$���@�,�?$���@�,�?	���!���5Z�H`ԒU |u6B����i����y|nI�U�V��PQ���M�I��
¡��*�:����8�А-���x�"l��@��L�	����OOVf�Xh�4����5��Rl��M���!#���'/�9^I�Y=��I�r��4�ׅ����W��~�
�#��*x	2[d�WR��x�Z��a9	�x�+��MHJw�j|�)$	��d��$2�[=7s��7i�2��Q�Kf|<ط�	[Q�䑁�F���$K` �C#���%�32rp�������Ty��0�uU�*䶃��U!qr#�0��1�
�C(c`��1����o�{~c��A�3�1�`*U����}~�c�f;c�f;c�f;c�f;c�f;c�=��)�b��)�O�9? ����f9c�f9c�f9c�k�k�dNa�-�A82
 * -0�t���Ƙ$�'��O{T����앰�y����}A��S�u:@�N�S����n�i��y,yq�$q"ڗI��(�ʃ�W���Q���+�C����&���/^ ��ŋ�7�|�#u'Kbr؅|�_>���5��Nm*&�А?n! ��զ#I��׍0b��B�ri]kaD��Qx�/I���.���pQ��8[��@hZ��M�b��>p�δ���z�}M��`��G��аl�f�v�l"\DM�|PF�_��׉����
8Z���<�l�������(q���a���V�;�T���zJ0^������T����P�l9"m�Dm�(���Sc�k��:�%�քk�i�ZD�^���
�%�8��Mz�#M��o'r0���*+J��kUz�Lq������5�u�Q�I�L��u6[JA�,��:��$��ܿ���֦vV���gc��x�r��H�u�y���)h��^!,�]q����q��1`P*!��F���&PD�t�Zim�Q PI$�����4\H)ڒ��8<I�g�t'.l?1�B"����0��N!|)��� �k��Q5�H7/m�k`�^D��b�Z�I�S�-�e���H�����Hа5�x�nVn�2� �H�UΠwR��R����&�|+Tw�Ć�q+��g��im�Hh'�A�%�L�55�#I�R%��D���W4��#�H֑Y����M��d� ap�x4�iM�k	�VjSR�	�[-��Sm�$�I��Ȝ�?;�&վm �٥,�4����4��q1��;l�,������}^��4|4m���&�6��@-	$"�.0��	�9< |W�ۑ��̸�k.ԛw�ҥ�)^��W�ҥsm.$�Ĝ48����xеN�&��96����i�&�A�o�#`,�6��u ��a5d&�l��M����Q6Bj&�MD�|�G���7�Ij�|��C�0:�L(���Dn87��H`�]MW�X�	���ƛ�lM0�0:�L������0:�L��������Q7B�&�YD�(��et,�n��M�걺V7@�����MV��>+�B���+!�stX�08D�
��"�0,�?/
��Y��5C�q�� �MQ���i΢Ы�x�F��"�먈F�/��㬨<����Pq�j���m�X����l,�jJ�3��7Q6�	c��4p�mʆ�[��+�[��bcޛn��ѡ�����6�b4ZZ��$kiI���p|�F��3����5�TlD%u��@֙Ԧ7V���|�O'QYAH�N�\m�X��֎� �b:'�y���Փ� ���h>i	��$Ӳ��sUn�v�>Ӟ�o���'��*
�Ty�'ߟ�9G3v}h򦍔M�%D�*&��4%@P�
�C(c`���� A� A�s ����9=�*U����}~�c�f;c������}~��__�����=��s�1Ls�'���r� �r� �r� �rr[ ��� ���i��ov���n��`��	�K��.O�M�
n�"l]��)
�6���d���������yR+%�Hc���W�R�"��?Q���#�l:�{+����b�|�~+���F^����� U|�I����c�X<�u (�#�|�N�J�.�8-S�nǡ|�#V=�o�s��|�!W +�׀�B���x��Ra���:�P
���5�s�����u�8� W����?�2ka���υ 1DV
M��T���|������#u��^	����x4��ȅ��<[#�cM�l��֛�Z�k���s�1��Lw+O�φ�mZn�|/U�I�iC��D�>�ς$ڴ��T�F��鷁�m�n�x��-WsŪ��8���7[U��>w?�-s�9�F'5��1{�<&�[|�D����F�0(�a���>Z���!���)>����J<8I��<�ߢ2�t�b�8+��Ԕg�U��7�s�>iBV�^/��4�HYR<��Ȋ��O��H�
��՚ɦ+B��H �kE���Q��#�"�kǓ݆ qR�Ui�X�$ğ�X�o�n�Ҍ�6��7	�.���Ȅڦ�ar�,�Er�ͪZD�pPH�u/���*��"nVjUr�ļF#B1��5a�$�H$\/r�\�x���Ć�_>f�����5�-#n�H���ܘ�AsSzL;�DD��؜S5�I��]jۓ�-�I�\�SBS�ěĠ��h~. DS�[�@9\��+\@@u��Ēr��%O��&�� �I�Sw��#]Ju���YvH��Gu��;���4������y�����p|�0"�jA�im*�?k���bE֡�#~��3R����Ҟ���I��b!���8����g�h~���9��|�.4,�6���ۆ)^��W�`�.,�łظ�N+cCx�ԚGf��9�Ű"�=�o&�A�o�#`,�6�#`:�i�R0�A�H4é�u ��`D�`~�7W�"�����C�D|Q(�椐j�	��`�:�ê�𚹲u6%���l�M����Q7B�&�YD�(��et,�n�]I��R`uԘu&]I��R`uԘV7C�ƘY\�m*�����F�C��V&U�Ѓ���$aa�1xT_	��F7Q�Ux&#_	��S���Z,^���a����
����3 "A0 �(d�ԁ��Xn/u�Bn��1�P�܄n����$���q�-�u~�N|�F��� ��	�Gc���D�WĂ��ݩ��kBh`��_�浰���,�>m-�e�����n�-8��J�����ڒ��:�DoMj:�ՀgZ̴m����@0�4$
���0�>	���M�Q�$[Wg�J�Q�F��&�'�A��RFĦ%Q����iV�+���xhL5;����ܵ>Z�?r��^�Q����9^�}��9Q�R��O�Ȩ�h\x�#�e�˙��C(c`��1����@
�{~c���������)����)����)����)����)����)����)����)����vG�#��1�S�1��'�Q���{���������5�Ul���˳o���ݰ
�*�Lva����;O���Q79@)��&/�(��KCA�h5���Sw��?|�&���i�	���NjKT�j�iބ�'�D F�#u

��ª��Ua���ȍ\e�V	��n�AgP`#� M�F�./W
��d���D��+���h��Ãx�Ԛ@O���&�uC��
��<�V8@?�0O�@0~�GW��A�&�=�O��d��3J�G/��a5���RvV���1Yx�+�হ�B�}I��R�ЮP8\���7s���I�o� ��A��)�+�<(�[i^)�G�{\�P<�`|�l8�-֕��w<��T(�7
<LW����|ҼSoƹ��w<[�a��l5δ���X�}+���5��nAs�M�( �~
�ªǷ�"�)�]I�EM��젼1>��-1��5���5'N�:u��/�Ã�:���ߡ��X���E��A�6�pPB�4�+px���zH����,���҂EPU!;�N��N��i6��V8�
H<�$ă�4>I��B��#�P)��2�yF^;�e��kBo����"Y�s�F����LY��G��aɄ#�M�J'��D�zԘL5��Ĥ����^<�G��u�C���F��??���x��N�+ᩫ���x�^�O���!�U�3A	�mX��I"��dR;��rkjW�k0j��m+~D��m�#�WѴ'�s+)O�YZp��d5s�Ҥ�vJ�4���Y��$Z�3�tqoZ��I�R��K�1$PSX���q��N��@Җ��-���Wֹ�q�ŁF�X� #�����7�B�`�%�J�$�Q@R`�MP�"2Z������ppm�1���ฦR��֫j2��\X-��T�qĜ.$V�ū�Ri�f��FZ�(��"�<�O-S�&�A�o&�@&�l��M����Q6Bj&�MD�	��/�����S��RW�D|H���`�LF���:�����uX��a�cL:�n�U��걺V7C���uX����ct:�n��Ɂ5r`M\�W&�Ɂ5r`M\�W&�gÃx��
រպjJ�7Αi����^5B��q��F�(���⠪��������0���<�*/�E����x�^5B��pb�� �-+Dj����#_7Bj�����*�n������&�7:�B΢��j�zG�5�io�Ũ���F��AԁS�R��%@�PԖ���AFo F���[���?Q�G�I �jI�Ri�H`�4�I�0DcB������������&�7z��B���W���hТ#D�������'��L�]0���Z<0�jv:�g����4+���Ĵ8Q�CjIX�REV���N�F�X� -P�~�G3sP��I���"��� }.������v�ٚ��`��1��0P�
������@
��1����v�`�}��L}��L}��L}��L}��L}��L}��L}��LvG�#ݑ�b��)�b���������{����������rOi����.A�@-�d�k���J�j��%Kr7(�$ok���!��JpVm��MG:��aÉ�7����hZ�6���� o ZG��H)�i�AAV�PU�i��i�B��Т2�4�_&�+��%$�	@�!�#Hq�i�V�����B��.jM��D_�_�����"�87��H��(��G�
&�b@�1 y�uzF��@�1\�W
jKR�Mfq�̾I��x��(�����*M^�._+�>u�cp�$���-|�F�c��x0|��:���Юs$��`�U㛹x�Һ��0���(�s
?��`���(�v
?݇�!���|�Ni^)�+�A��4���Q�~���У��ҿ�������<\�ηֹ���F9��M+��<� V?=�ADbp���^=��S��r�>nUOa7S`;=�N�u"��8�h%`��酏��F����hW�X\aV��6��j�d[E������V�\G`�,�ޝ���K�~ג#G��'"�=�� d�0� ���૭N#^/ޅp���/_�c����>^D�O�j�OG�N��u�p�z���D�u�A������i�e�U��&�u<v�c�Sۧmۖ�"JmU*���%-����O������qŸ>v�91�����x�K�S�"CxU�����(�u�_)I�"�|x:�J�������c$�/��L�i��R��x �00R���7(�*.�v[k^N��H���F���V,��"�h���A���L+C���鴂gZD�~Q,��v�9H$���V�|�=@Q�F:�-��n-L�1��c��S����/�p-6�0�P�6,��+I��Jr@�xq5�;n��M^�r qS#�&�����RY�|���%�ڌ�{Q�B��l\R���q"�4-]�f��Fo����j�Z����x��7��x�i5d&�l��M����Q6Bj&�MD�$�T>H��M#T �7:��4����&	�Ң7m.�೩0:�i�
��Ьi���uX�	��j����0&�L	��j����0&�Lz��B���_����|~�/�ޅ��о?	��!��TqR���<?i�J���(��k���F�j�׆�5�hAxZ#_�WšU�h1|P_	��aUayXP_�����x�I����P����0+�j����#_7Bk����*�l��͑��&�7+j� ���|�-��j"��HD�:���"ЃH|V(�"��D`W����U�W��gR`YԘuMP"@��7$�J@����J��,�-	��a��\|V���5�kЮ-+��ā~�F���7�I�֔M�N�cf���n���%�U�I�?��J2����K���Vz��-~��jPo	�jq5��.h�����Z��Jøf�k(m*ִ�jl���U<z�^��l��$ (c`��1��0P�G�G�G� * U����}~�`$x$x$x$x$x$x$x${�>�c�>�c�>�c�>�c�=��)�b���r� �r�aWaW7���������n��D�}D�	r�%���kh�ܥ���Na4�N��ĹhB8u����r1��551�~�G@� )FHQ�Ī3x��7�����#xx�-R��%�!�7��D�Y"\�.�-N(�S�C�PБ\ԜK��E"�kQ���k$a6�i#B�.8����͡��"]�R�"�Ґb���ZF=�'��Di>I�(���F���Y���M�<�7������x��H4��
�uD����0���.�:���r~Ԓ)�B��*�_
zAA6��:�=��A�
�p��`�|B� /_=�׀����z� �&^�/I���Rob�؅x(�}
$�71
MlX�[8VŎ!{��^�{
:��b���CHǡ�cТDWcĚ8�X0&�8�ۘ|�ڒ��&� V'��W!�,bA�D�,�V��qo��_�9`�>ky��ƹ�a`#�k�a6�*
B��̛�W�hZ���V::�����Z$F�"j� .����6)�m�� �:���tF�:ǂ
�1zL�^�0����)�|�Y7��4uU��#�x�ГpI��m�3�4�ɊG	�j�#Ua�H,^N��Cn!`�:Ԟ�~�l�܀=��ShD�l(�[��,���];����B�"�[��rX��6��a{X�4�@�?�� !	��E~4>v�-���|��Z:�m�_��д��p���1�g���IM�hƁxXX��_��M��nnGQ���ޮ�-1���2H�u�)Υ��$��|btuC�k|i�E�u�Q!�|�j�5�h|�yJU�-$Pw_���w
�`�Y������Eb�D��|�����Lh�U+Hl6O[��;>ML"��Ѝ�,�3�z��BG1�`�ph����8��:��Fm�>JQAe��JFq;��qJ�.8�����БsQ��7ɼv7�o�H��4�ϓH�H'��	�d�xuD�Q(TJ��uD�Q(TJ���l�������RP���u��Gϓx~ԛ����n�+��j�����_4�
��AX�V&��sd �l�͐���W6B
��A\�/���b�0�L/���b�0 �>|��x9 Т#y�NGQ=0hV	�c�3��F�*�M�nq��F�78M�ę���7
����b�L�#
�
�⠪���>
��«ƨUxn_5A��1||#^6^��d,�>	���k��U|�z��5q�YX`V5��%�u��F��1DDi	�����4�Ij~Vׅ�5q�YԘW���5q�M\nV�E�gQh�Pu(��5\TV=
�Ђ�� �0+��� ��� �"zh���W���~�u�_T�@�\�������x,�/�����c����?�Ǔ���Ks�R'w���ݸ��C���4���RFġn<�4N�����/� �AWÁXS[F��%���K�ܤג:��&(c`��1��0P�G�G�G�G� *U����}~�G�G�G�G�G�G�G�G��c�>�c�>�c�>�c�;#��1�S߮A���A��7���5�5lll8@e0܎�?[2�sT�}�;[��	������d�GR��?H�jJ#���e�4����"�RZ�m-��86�kQ��kQ��"Ƥ�cRZ��8�>JT��nq�m�(͹Ƥ�84,������Q�*IaQ�W��|�W�#8�2FԒ1q#����@qS �N��`�?q"��q��[iZ��(`�#�Ԗ��b��<4,�3b�����'�JD��<H�:�`Y�<H
zi9���<�&��52`~�Pm+ B4� ��,�8H�-Q�����@�MDxF�<#Q���E�����Qpc��1�\�8u:�U�B���U`��X)�V
+����������_
/�?��/��(�xxX�<�#�)B
�O�H�ɼD�V���*��jJT�!vґu�+�۩���a1�Q�B�?o��X�4��|4�8�-b�YF
GΜ\jA@�~jOL�|���-��?_
�04��S���EF�A���Q7�5N��)!�D�+ �����ۨ>M�xA�>/í!hUXP�(���sTpY�C�R�HF�]�'�x�J��x�M��kI��MI�HΥ1�H�=���0L���Y��M��x�n���dԚR
ebY�Ҿi��%�*��ĐI����c�|�(�m�|�x���:1���Å֭W$֎��������V,���D�H��!�J�'�)2�u+�m"���#�{Z���$�xa�'dtr�iNk;��H�oD�u��UP5H�7�V��L|�ECCH|�$��������������$DD��i�p����F����n�Q����x�c7���9^8^U;��|�w|uZ�xu��'�1ͼ6�xb8=�JT���Nm-��k.�)E֮�D��Б[I�BE�Ԓ)�2��,�9�� �A<,�O$����@:�P	��7S`&�l�M����u6n��M��	��gSe�7��2@�&�?
������c��&�?Q�F�M\nW��Ъ��_6B���U\~#W����`1x�^&����`1x�^&?����|�8O��	���>'����I����*��_(�u1���(ס&�+�i2���F�>�τn��c��X�?8O�� �L��W	��o�LF�*
��i6���>'�U�T*�7/����A&�zmв��,�?�"5�e�_����ea�M\nҼ�`�n��|Pu	�U�B����L	��B��k��$+JA1�V5Bj���D�z�W�|�z�W�|`W�U�O��M�V	����|Z�/�C��ס\ZV���ahMX`#I���cc�@�>H	�%�ڴ��ݸ��[�i�ï�7�|F#W�E�5hU\���@|$F8�H&4$ǔg��\^>u�����'��	������n+Q��� �H���b�1�ӑ�W����j�{6�A�$�#�~�S��C(c`��1���������A
��__�����������������)����)����)����)�o�7���3�1llllllm�
�
��� H4ߑ�T���}\�}a���><ݝĤ���sB�ܜ���.7�q#jKXа���(��ͼ>5�d��$mI�1q�Q�a�C���p5�ƶ��f�?Y��j���|۠)X86��Ұ���X[K�4,-I�P�JǦ�ޚ� �D���~����
X�۰hm�Ԗ�Km+M�`pp5���](|�.46�g��ajK8��T��@���X5~5ԭ�&�kl��J�Z���C9��\XGJE��DZ����&���"	���⠃x� �*7��"��H� �.��F�H�iC�Ɛ�U \F�.u����G���@�R c�1X����b�P�\��H*� ��VґJ.)O涀"E��	4��<���Ē����J��Q{�����Z<^s�ţp��N���/������j&�?�)yٯ$ 7~ �-0_�(�l.�OK#fA���p��!�Ұ?)T�"xyD�zFʌ�n���MD`io�0>5�_:�$�({2��B��G����"Ab�����ט��@��	504����datqH2e�S��MG3��]i�=��ko��˗v	�������0`A���_S�]��>�G��	8��ǒ��Gs� ��uJ�Ҟ�(���<�)��S@��
��u�N(4�m���X#�.�h������H��ַ�"a4��-~�I�v��;�J���u�B����:�7Q�B0#�ڳ,��\��\ԤR�B!Ԝ b�jBд53�*���ځ�X<����5Ͳm�Å~ԛA�B�&ŧp��V��ք���v?�m���OjJP@E��M"�i_%��io�J�A�-Zj3x�|����NzE��D��(���A��:�S`F�i�Ս0���u6��A��:�S` �l�M�"A�u&͑b�0^�L��5���&=�м>$ۯ�M�,^7E���b���+��U�T*�?
��©3�L�*�?
��©3���|�8O��	���>'����p�?���Tx���צkj����pܕU�`�	 �&Tp���g�7Y�1�|p�'���Q��
8L�2������
k�ЂM�p�'��	��&��ڢ4��A&�zm�����^?�����l���B��:�-z���T|�7�J��� ����/
����b���1�N��k_Ǌ5��n�1z0��_5Di6��&��ڡ�M|TW��Aeq�-|�ů���:�-��^�aSЬ*z�@D��о#���e`�RW	��$ŹO4����ܨ��ϒ���_��d�P�Y�0-K_Ę�YD&#p�?�����Q��m�|P�+��ħ�uZ�jkw��L��db��p�Cβ&��DZ��`��n����6����������j�.��Κ1��0P�
�C(c#�#߆_�C#�#����A
�{{{{{{{{}��L}��L}��L}��Ls~��\�1�3�V�V�V�S�؜���T��'��=���6�j��j�hL?~��۳Q$�HO�3@��ۙ�*���-b��.$c��.)cB�4,-I�jN+RqZ�F.)b�)a���{�m����u�;r�ΦD��ȃ��~ܰ?nX������l�qqg{RY�fޣ6���
[�Y���4,>sZL���ͺP��`~���X~��v���w�ܱ�,p�g���)��v.?O=3A��ۿ���"������Z5�1�`�����T�Lֻ6���\H��Z�+@Ц88�����~�<4,P��qF��\Z�$��$�$�R,�XH�:�`Mj�Mj�M"��Z�z-BE� �JZ�7��"��A �A���$&�Bm�_���sjJT�*��������L.��LGF�B�xBu�E����B��k`��E�F��>@A�� �(��8Q��Ԅ`G�@һ��@��Cy��2iz��`���=�m[�2#���h+�M��ք�J��͉�B�8,�[7��*��!V(�*��<\q�����U ����A��({2��S��bH&�kU�r���6U�ԬnI�W7���%MQ*�9���Uh=�
.~�PF����#F�N;Tܠ��$�I,�Mj�d׬V'E"���I,�ė�%����S�I �������tƛu���:S��Ɔ \���%˴%=D���Q�;M9l��й8Q�6�szH&$�NnLGua\��d��J��IFQ<�K�M�u	R��Q��*����E��&����ۭ��H�R)�N�%:��Z���b�4���� �X-���#gI�w+�h1ۈ�Ju����ӷ�����j�jk23��͎m�ĶV'�NOCH�H'�#H�Q�F�u �z0b��u(M����u6jƘ�X�+� �sd�l�͐b��W6A���1\�+� �sd �l�J��Y\�
��"�`�x�,W7Dj$����#I�Di3��M0^�n�Ri����|n/_�f����p�?����|�8O��	���>:ڡ�[T<�j��mP�u�Cζ���|�-/�j‛���eJ�fTu�#aT�@U�`u�fWY�y�`p��f+��ҿڡD�hyx&^ׅ4�P��nu��g��	�1�n#I�Di3���1�I�^���Ax�,I�E�6�1x�_5^��оj�M��x�/��j�𳨴 �:ʂ�ƨAXZ�6�#�:��c��\Z��i3w��PV7B�3�L�*�?�ڡ�hM|TW��5�hM&n^���A5�PM\PW��@D�hY�P#I���Aԙ@1��jJ#��,��Wc�gQh�&F!xRda7Qk��#:Ѣ5qPA|T_��A���"�7	@u�D�+F�'� ��($Ȃ���`�Q�6#V���1�DZ	���t&�m.�0��x*Jz��C(c`��1�����/�/�!��h�B��A
����c��=�c��=�c��=�c�O��>�D�)�O��>�D�)�A�������
�
�����'��=��lPsca����k�S�F�n��vhS�f%J85(�l<��>u* �J�~����H�ƁiJ��R��tJ�f����q��`��c�5�9���w�k��~k�F�~k���>SC�4?na�sۘ~�����0�����>SC�4>SC�4>S_;rǦv��4>Y�͈��鄑�wΦ\�ۖ>u������,�ǃ�cB�SC��8�����:ɇ�i������,ۘ��2u�[�S���ͷ4�Σ[ظ�<Y�F+��i��e��ޚ�p���N(uK,!�F�mI�|��a|��a|�W��|�P�FH��(u"�� � ��PMĨ&�DH�Z�[Б�	uk8�d�'��8H���N�cA5�D1���
��w
�7Z�
5%z>��q�ޘ0>|��W��Z��lX5ݬk��T ���P�P^��Z0�ژ�%Bk�3h����-7v8��U�srY jO�hMڇ���ܭ���E�pYJ�#X9�\O��а{Q��b╦�ԧ�3H`Z���7ΦP|�'�|&b*�S����Ij�I�pꎓn/�Ȍ������\z�J�͖���@0���-@�!ra�ࣾO�Qz�+�J�m��,���&�,K�[�j%}m�g�7�|5��M��𽿽7p�������7Σ��������C��$1Ɍ�x�K`\�v;���d�6*T�Lݪ)�"��@;���6��LR�����G\�S[��V8J�V8
'�J�iUĂ����6���Di�`�'Ӗ�N����Sm��&ܞ6��bY,�S)��!ŤiGbz�DL;��r`�$S,��D�srvx��"�|�_�ہ\��Z��ct*�P
���Ű��<,�l�Mг���Q�I��R`yX�
��b5cLF�i�͐b��W6B���U|�
���U�t*�n�W�Ъ��_7B���|���5�`X�l�Rm���0^�LG�C�0�78O�����0(�?
$ς��
��^�j�������y�|�������y�|�:���Y���?g����u�����c�1܌l��b�	���H�$�f��*�$+
��Ы��*�0
�KC�2���L(�$�So�����p���eU���xP�$ʞ�	�A�`�A�pc���>�S��A����©3�
M�!p���4�M�^���B���/�4��M|~�/�^�X���*8O�� ��L*�z�����Q7BΦ��P
����4��M0*�?���К��&�*$ڡ	�A&�/�⠂�� �(+�
′@�F�(�OB��u�f
3H�Q�#�W	YX`u���ס�`#��U�b�aP��Pp���P�ČX� <F�ǀ��n�
&ȍ�&##Q��
2��F�?ǃ���xH^��"`�q0�0�>u'�Q�c��ݴ�
�oh��
�C(c`��1����/�/�!��c/h�H�H�ї��}.���}.Ǳ�{Ǳ�}��R'�H�E"}��R'�H�E1�5��m��[{��>�j�˳.t�i����7[�9]�Y��ho��c!�8pۿ5&�P~�Ɔ݃C���~۠�?�ƵA�nx8Y�&�C���I��O��h���v叜�|����ѭ�ѭ�ѭ��r�iM��~���5_���s|�k�6E��靣���������h�zghpv@'�q+�W����й��#�]�k.��ʕ�� ����]_��L؉�ҽ3�A�W�'k�+���r:К��b���hX"J����l.�
��-yv������鍡J>X.m'h��B%OL�e��=5�!q�)af��[z�XU��4)m������[{im�Km-���o���)o��X0,�DR��V�%OC��ă��`Y�8�gFXZ��ԛuÃr�8'��OcCxF�m��u�!b��A�@?zb0�\k��WHX�癿�گK9?�`<.@Gp��]%zu����R�͗�L��$ 5;ޢMT��a�QO2]
H�8��ɠ�����Ă{�܊��`ċ�Хm��� B4��Y��ԖcB��o���u�?��� �MGE\țe�"m#�RAbSxԞw��$�v8x�޷�4l<1�rz�������b���hn-ũ53�:a�E�a�	bM�f|�X�^F�*��gW�߀[�������2?���,pX���`���-�U�?�߀��~F�m���-����p@�;�64��@�j��q��80*����4��i%�_4�*0�y�&1�/�A�����H칞\u�u�n�l��� k!�7�G���f�|��&ҵ/��r�Ɠk��N��F5X�F��˽�����j�)T�㹵A����v21�`�*�T��W2�G<���4Ɖ,���baW���0-_B	`���W(=
ƘuԘu5Bn��UX|,V��Ы��#V4����1\�
���U�t*�n�W���x��/��c��L����1�^&?���u\�	��M�!u�)���t�l���y��?υ�����>u���g�G	�Q�`/u�C���{��^�>
?���{��^�>'��	�1�np���3w��|,p��]m�{�m�I�4���
0��V]cb� j�p���&�	hy�Z^	���AE��xP��8���YhUx&I��bb4�P��nu�]f���p�?��𫅺#u�B��&~I�\-1��I��g��T �j�m����*�>���3w��T�<��h6ib��l�-+Q�4�T,�l���L�<�?$�©3��#_��A5�h�&����i3�M�^����PA|Tp�>J#����<�(	��j�Ƚ�n!x�eC�4*�(z�7X�M&n�+�� ���W6� �^�d@Ę���7|��P��_������V����cB��,�Da����������^4�`�cB��Fp����0��s1��0�� (b�0a��4r�r�������2�^�^�^�^�2�2�vG�������G�{~c��_�`.@���6'� ����j{��j�0MAr5��5>H�N�`�"����Gc-L�d�64�f�if��7��ޛszm�qnc���L��ܠu��u��u��u��u��c��?-/����l���c�c�c�c�c�d�6^�������:͑h����蚙�������
��v��i�O����]q�W<u���s��=�+��m���	����5B�͡���7�榦`�ܴ+�h�D�&���&[���<��lQ��
u����B�j��[�Ozs��	�,���Ƥ�T-�L�ǟ:�pp�ť4\Y�e���ܱ���o|��ܰpnX87,��pnX871p��ѡL��LƤܠԛ��r�RnPQ��f����m-�hRƅ-�8��46�BL���ɋn��k���`��?��Pz ����ɱTF5  ���%~P�:����z�͡��*Cv�Lx���_�C��6�M=��$��D�V�����f1��p�Kx�Q Q�����1`�F�.�Va��X&ҳ{�A@��#n,�i��� #H�:���Hޝ�ݞОE d�I�z�7�H/|����׽�l1�M"���b�s�ۓ�tq���$��;J�,��m��~j�X��0X����>dW���~��di�l��o���_������%�?���߁��~F���37�o�o�������*�7�o�e^{�g�7���zBگU���sXߩ��i8ת�&#^���N�����[�k~4�l4���(��. �8Ǒ�{B~2T�F�������%J��chZ��i3�A\�z�'���GY�X�#�0rrDD�>n�%D��Ǐ\�URaXԮq6��NI�C��� 3�BT��a��<�*�*hTyq���6%w �΢_�W��D�M�V6n���|�,_4«�ȍ\~�+���1|�������x�/���tX�n���b�,^7E���&�/I��i���`�&�/I��i��`A|�m+Wg��~p�C���|Q'������u�?��ȱ��?�"�Z`�֘,p������Y�Q�~�:��nˍ��i]m�zM0&�l�(Ы�lF�#�F��4(�??ۢ7[L �i�Rg�Uḍ|Z^���5ḽ|n^�&�	hU�ZI��b�qk��i��¡����C�0��� �?
���WYC��L/��T|�l��m����_4ޅ�dF�i�׍1�#^4ޅ�e�_7^��tF�L�S	6�ГLz��5��оn���\~#W����B��F�?���j����F�?���j��b���j��Q��F�7�ڢ4���&~#I���mQM�#I�Di6�Ax|^����Ax�^&���`A|�/���T �j��оj��м>z��B���_����\|�+���a�M\n�/
��CГ*zeAԙPu&TI�>I2�|Z_� E�S�(�ʃ�2����F^(��x`�/�as�.f0�b8�@P��3G/G/1��00�=��/^�2�2�2�*�vvvs~��__������-���4�'�ӟi϶ó+l7ND`�*N�����
h�S \�S�)�`l8nQK5C�Y�?��LָqS 8��T�*d2���L��ܠ�M��n&�q6[���M���zgh~W��{�;G��6G�靣�����v���zįn%{�'���H�𺣨$�rh\C+�8'��D+ڙ^�	����hD�	ꎣA��Ohja&��\8�������J�Tț���O�Ge�м"\?���b#�4��9���̔�Iq�4�.y�b���8LG"!J�Av�2c��d�)�8��E)�γ`⦇�~���eO�L�Z6^�sW�h~l@?6 �͈���b��v`|l@>6 Ȇ�2!�L��7+�I�si6"m&�MH��qgx఍�k�����-)S�Mx���t�#�����$H:ֺ�ֽ�'M�V��'�B"�L�b1�&�i4��LM���@�y����bc�{�9�'�맙�b	��I�c���p��@�j�u�]�m�G�n$�If>5��7��`�H�,^��`:����*iXy��t�C�D�S��Ÿ:��"ˑL3S^����e��#�	v����ڭ�4�6˚���b�zj�
���,v4ȶ�K��y�4��F��*�Ŵi����Ҽ��7�o�h����a^Al7�,y��cϙ��4X��r�h���n����O�>f|�X���<X���<�y���M��������|,

�^�%�?�l�­�q_ 06�m�;)GZ���S����%�n5n�=bT�(Nw��Q�=�l
A�-I��4^�6�^*@�����Z��1�
����1`o���<��O2\�ʃ��4t�1r��w�O�2p��*��#����� QH��b�Dcd�R_:�� UX|��/^	���xQ&�/����A|��«ƨ�x��ŋ��x�/���tX�n���b�,^7E�4�zM0^�L���4�zM0^�L�����iZ�?���1�u��'�e���Li��1�u�?�����l������l�������<�>:Ϛ�Y�m��M��c�L^�L���г�����c�X�Q|��![t&�L
����ƨUxn#^���4�T^�>�3�{��u��fU�h�X`�+��\T����L�(:�Ŋ�����u�������i�d:�i���Гi�	6�Гi�	6�мl���мl�mЂM�I�^��u�_7Bj��M\�	��!sd �l�͐���V&��b`AX�V&��a��\|#W�Pb��_���`Ax|^&���`Ax|^&=���|�z��B���/�ޅ�u�_������ �j��P���_5B�A|�/��B���W=
��\|�+���q�Ю>z��5a�YX`V���Eq�\nW���Eq���0Q��
2���*/
����&P�/�%��0+�˙�3.f0�˰P�`��G/G/~/~/�� * TP�
�H���\߮A�������  �ݰ���S����r74/�6_P?vDZ�M9j�yB�n�FI$����c��j9�k.-)R�JT��r��'Πm��㉭Q�va�va�va�va�va�va�va�vcS+ڙ^�J��W�����9^?&8Jc��1>�	��n$������-�����n$�����8����C��!ɢc��9��
�)^�	��O��|
D���DI[��+h!4�ցh�q靚�^^p����L!%y�)T�y�d�L&6��f�v8����*L���K2�4�Vn��QI��Y<"�����Nu��L���<?��Y�c�/L��º���zez�;1_�����W�f+��ُ����v`~W��{�;1�8�.�����p؀����೎8���e�pSC�}�$k�H��K��Uk�� e�RUȕj��a�J�e����ޯĖ@cc��5���전�+�٢N N~~+��#ϒA�&�G|���f�`1`1�Xm-��f��6��%+���v	�\�i��?(��
�1��n./��p&�Ƅ�%Q�k����O{-��'7�&#y��ʘ��Z�	��ѡ������4��RM_�b��X6�zX:B�b��X������>|�X�c���؍0-�~"���ߖ?"ؿ�,r߅��c��/����|�4�~�_���et4��uy��?�,v-�Mb-��ň?��������_�?�����Ӿa�(����mz��n�N�ٿF��,K�zE���g�XR&����c����i�N�+@cqW<���H�T�P�7շ744�ԭ�DR�JBǁ��󘞇���6�F��V���Ғ�D��\�"J�q���]�����ò�p��';>�E2\��LD�\�@'�H��D|�d�۩�A~�+������n�j��0���|�i��i���T*�7
���ƨ�|�
$υ�4�zM0^�L���4�zM0^�L���4�zM0^�L���4�zM0^�L������r�ڡ����|!�C�"ر�~,p��'��	��֘,u�i��Zc��L
�ς�����(�Lq�[-rM�!I�C�4�����p���Q7�ۛ��b��\�+� �Y�1�|!I��Rf���1&`#p��&��st^�n�Ri��`�&~#I��������V&?�3q�?T��"��*�-+�Ŋ���D�(���Q���l���xM|�	�!5�L �i��0���_4�
��A\�+�"5�t �l�͐��1�u7^�Su�u7^�cM�V4ޅsa�W6�sa�V4ޅcM�V4ޅcM�V4އSu�u7^�St �L+
����&�L	��j��0&�?	��j��0&�?	��j��0&�?	��j��0&�L	��j����0&�L	��j����0&�L	��j����0&�L	��j������H>I� |�(��e���n�Φ�RV6Teq���?Q���E��\nW����|Z�/��ƨY||_3.f\�av#�`��
�C�^�^�^c#�
�~)��~~``��� ���d�
�n�ۯ��&&>��}A��l�Ϝ�9.*[TF���Ʉw���-���z��҃����WT��*���p��Dc�jf���@�q+�Z��W�����įn%{q+ۉ^�J��1��h�f��h�f��Oa�h�A{p���:����$(�"�B��6�DS�1����2_���
�DP�6�`���!(D%m�h	@�y(���Ir��xrL8'y�k�@��B<c��I��J��&_�я�s�Y$��j7x7'�3r��1�Bb��]DVGm��M�}_6��$'6��<�&!���JV�N���z1
�M�W�a(�"��uÁ<��WA鄯L�zf��4^�����h��E_�*��W�~W��x|W�fffƆfh�v��h|����.70#o��E�`%du;b�*Ta�˕"\���˕"D��d�'�'�2�(ʜu�I�� �|1s6hhW2yR� �� K�!��p�>M  ��3аR�z���J��6��%+��v|�I�D�M�o����<�7����Y���mJ�V�f������;�ͪ��d��5"R��%7"�*�<������nI��sx"�n[�@?k�4�W���X�l�����ߑ����r�e��c�y��[�>|������o�-��� 4�c���ݟ2?�n��~y�M7�W�4�b���e���_�,E��/���|���^G̯��|X�����W�xi_U���|W�����,K�k~1n-���-���/�o�^Ah�&���������{�<??��L��55�0"�Y��h���v�G.0l?7�\F�	_�&����s���5��ӹhV	�M�	d��vT�*%HꌗT��1�ChPOl��D#K|��B�a��G\(RU˫�\��%��Ih5:���&�+��γ���ҸS���&���
:υ�3w�&`,^Rf�*��|�?���4�zM0^�L���4�zM0^�L���4�zM0^�L���4�zM0^�L�����^�j��g������7�a�`y&�I��i��`y��8[��t*�L:��i3��M0^�L
/!D�`X�l�mס�`p���צk>	�����7�X�
�����L�B�j�W�P���F�7$ڢ4��UX�+���L*�i�	6�мl����U�����q�~�i��g'�D~�$�����yԘZ��A�M�l��UrpYX��/��B���+�B���+�B���+oB���+oB���+a5d&�l�R0�A�H4é�uԞu'�]I��RxuԞu'�TJ��uD�Q(TJ��MD�	��C���:��et,�n��Mв��Q7B�&�YD�(��et,�n��Mв��Q7B�&�YD�(��gSd,�l��M����u6BΦ�Y��:�!gSd,�l��M����u6BΦ�Y��:� D�` �H&6�e���-�D�m*&�iu(6�M�+-IX�jN��iV&6�Q�iu(�ƫ�?|�ɏ����W&3f0����`a�1��!����������o�~~b8hg���*��@�
~�?v��ϟX����dM�e��dM�T���)k��z�*C�^o'�L�D�1�˝Fĭ��cpSN�e���1�S%m �hڙ=��Ё���)���)���)���+h�@6�����`���0��o8�C�a{�"�����Ju��1�"���8��S�	��R��)�"� �����EnxDn&<��&#	�#	j�����,��KJ�
m9fu�m�D2b��L"�{H�
�s�Иj�����iA�����'*��+�ϪS�	4xD������P�2�z����'%��RdZS4e�9.�������ǦBT8��uC�6㉢��>��>��>��~h��D?+��?+����?+���/�����M����6�x|kGnw��Hx�6e��^�UփȚhJ�)�/����
 �1������z
�Z�H����e���]�<zƃ�E7\�7���p��G0���*�v6�A����}|�O�g�u"�H�(��RZ�_&���H	�F�*LM��M�oɥ~~��e1���#KW�DǓT>x���m.�[JC��"�L�&��"��*y�BxTZ+��DYo�o��@�jϓ����b�����j�|�<�B�O�5|W����,K~���+�|����;�/�E�|X�c�l�݋�^c�%�?�|X���b��?�,D�ض
���_�e^x�E������0Ӎ;�J����W��c<�B�?�Ѐ0|�iZ��'���p���E�%�6�d��8u�u��FRM�~�'��ώ2q����+��B��V��͠.�n�ڵ�q�����Kz ՙ1�n�9�.2����☎��;�+�cM�JI�g��4�Ls=�v~Am̻T�8a�ʙ<�e-�:��A�P�L�:�j��g�+��>I���kn7�u��-QzL��^���T|�j�����`�&�/I��i���`�&�/I��i���tX�n���b�,^7E���x�/�U�u�H�f�����_�g�D��U|�
���U�t*�l�W͐���_6B��ȍx�$ۯB�#^6C�����l?���1|���C��&��B�i�>|�E@��P�X�̀���W7D*��
��*�>z��5��оn�
$�b�<F�Nz��e�pY|�u(�
�u�V��V�p�sQ�E b��Q'�]M���n�ׄ�5@��O��oC�9���A5�L:�PzJB�A�Q(=
%�D��(���Аi��F�M�l�F�uj��[ի`:�(>I�� ��$�$���r|�O�Am�H-�I�� ��$�$��Y �Q'�	�����((��aFo
3x�Q���6f�7��#H�4�0#H�4�0#H�4�0#H�4�0"A�H'�	�D�x �H'�	�D�x �H'�	�D�x �H'�	�D�a�Q4�$�e�H6@�&�D�:� �� #�=�����pАNjI�RH6J���TM�Ңi�Φ��l>N���l3f0���P��� T<=�S_��_A_A\�S������n�����Lvcu�u�su����qRr�r�؛�ޡk�!wz��d�&bM2��Ɔ��W�3��;Lse��-�Ё�h\u��7z#%:�U�m{h�@^�����m��n+p[�
�V�B�2������BrB�JU�1���N�D����1�92����"R�D�q&Lr�![�
�������Rc�Ba(���$�<�&48Ik�cU�j�Q5�G'�E�sJ�j��'|�6�d�Q7� D�h���"vi������M�rB)��w��4ˬ��������)5N����iGx��AejbT�5_[q4 ?��+qC�D8�n$�C�I(~v~ۓ�8J8�#����>��>��>��~h��D?+���8������h�|���6C�4>SC�4\SF�d<�24�L���h��2�l�w0vh=b+ ƅTk��444T�t!�\�W�ӊS�#�JSX���UTe-r%ٕ�5��0Nrkʜť�����ZE�c��<�O$[5�xYj�Z��֫a�l&�6�#T�>J$hMD&,Q4��&��(#
gu�������c�h�bF���!�B��x�E�`�Zi>����4&��'�j����m'Y�;���6��p�������w�?����
9n&1�-7�.#�i|��t\��?���A�Q�`���B�0��:
(�0x&6���>w�zc�iG�qƁ�����Φ�8���V�G��c�� h�y�"������Pus@15!chZ����t-�)��(�TM*�ld�y(���o0��B��<�Ko�i�ʕhJ���03��� ��J���h�+��EWa�B�T��U2q�\���l��@Ux&!u���	��c\�l;����`>�E� ��I��������\���"��tX�n���b�,^7E���x�/���d<�l��͐���_6C���y|�/� �sd�[/��sd�L
����`�u6jƘ�X��5c`F�lՍ���#W(W���MX�V'���C�9�u'>N��"��x�(��7Α>$�j���ԜW'JU`^�l�����Q7TgSeFV6$��YD�V9�M�X��U��d�xu�P|���о0jM�c�m��e��Аr���BA�.8�¯�u\:��i�2��,�9��PAeb��r7�Af�l,�9�Ű�x�o����u�N���e�xYj��$S�$�s��O|��J3x�4��f���Q��e��7��3x�7��3x�7�j3x�i��#��[|�mIj�Ԗ��I"�Ԗ��I"�Ԗ��I"�Ԗ�ͥj��[��ҵPm-�{iZ�6��=��TKx��[Ŷ��-���m���m��[m-��io�Kx��4��3H��4��3H��4��3H��4��3H�H'�	�D�`�O$�er��NQ�KcCx�47�cCx�.4�b�H�.4�cCH�4$�ez��Om)�ҐNf(�Q��{�xdxdxd{����!PB��__�o�7�sݰ�l>��m7j����P}�>���a���&����CM����4��b�L������c��y�N<��6�{A�\����:�V������ML$��DcX��K�`k�r�����n+p![�
�V�B��&Tr�G)Tr��&N�d�&@���%$2d
K�]��9:C%�%�Q�Ȍbs�drR�
Q�J)L`��ۀ^ !*��%&�rU�4@DDL�&�^�<��d�A1�.У�gQH����DbT�64�M�"D��7��ƽ��i���E��DP�Y&�(���ķ�j�SI#��J�kKù�rhcY90.SPm��W����(E1�W�lTu���ШZ�jd��10��ܻK7�O`�h�xpW�{�4^�����h�Ex�W��{�;1����������-*�����؀�D8)�
fV�*$w�����L�HE��f�j~���6Q*h<\2��g��802�H����@�5��f;n�jJň��R�F�2\��˕Q#��
2�A9�"N�w@������x�-Sm#d,�6m#`&�6i b��Q��E7R4&�4�O���?R����~:��9�.j ?n
R���8�kAM�YM����b�M-���y�sk���Юn_��4��MH�jC���>v�#|���p6��
�D/CR�
3��5 �|�E��F�~:���u!��@1���?���4��>�|����\��oCJ	����\���҇�ms�
���8��qQ�@���4�N�R&���
k
M��F�4� �5�H��]�T��@6���)��<���2�X! P��
O���[|�OsT�Q�H�=�Pe�_��j��_���j�t�Q��i�� q�&UJ�!���z���n爚m�`�u���m��1�x�Ey�`I�W�����<�n��́z��W4��sM�W4��sM�W4��sM�W4��sL*�lU�����V6���UX�
�Uc`*�i����st�P(�Uca�,�="؍D�#u'�I�7Rp�Ԝ#u'�I�B��:�r:��n�0����H;TN���iH>���M�`p�	��n�Ű#x�#W>��Gס�s
�\�kU���=�7���H�4��I�[jM#�iH-�����Ԟ��
Ij��R-1qĜ�$ʃ����P|��g�jFX?(�"p|��+��lqnV�JEʹ�_C�+�ԶZ�����d��Yj�H��.�d��Y"�Z��V�aԋ�Y��q9��No���Fq>�����KH���Kx��Z@��{m-��RZ�jKP�j��[Ƕҵ}Q��e�vQ��1q��.8������vNB��\q9�'a�"�4$\Ƅ��Бs+cBE�hH��	6��rjM�Roړx�ԛ�6��9�&�ͩ7�m��rm-#�ii�KH��ZG&��96��ɴ��J3x�7�j2�ɩ7�mI�sjM#�Ri��H\Z����!qj�.-]����ho����hoƆ��hoƆ��Q��1Fo���!����c/c �A
�}~��\�SO�Sm��M������%�I��O���&ò�d�h��Z�(}�۶ԒOo�4�c��a���Q(Ey�����+S΢e��19����p)0
L�Iw��n)�DcQ��M��n+p![�
�V�B���Q2u R�"R��*�L����!��2t
K�j����KAND�'"Q�ǛA,�S& �	��K�%����	 (^���]�A'�H㬤e�R2�)#�A�f�r����F+�'�5�2Z
9I�9I��\�J�%�4,�[��f�X�
�k�]4��'���5��L��8Lk�֤�M!L=� ځ�p	Jm��aL�D.�wX�mN�jR`%���"l2L����hA������鄑�bYè��,�Å��W@~4C��8+Â��/L�zf��4E��Z+�9ُ����v`|l@>6 ���W�h~���h�D8)�
dMI�\.��ZH�
��
'��L�u�\F%��61�480R�ǎG2��~SS	�. �Ե�Y�͹i5�]	s�O4%U\+ޔ0ǲ&����=�RBǃ�Fu7B
��U�>4�PbA�Q6Bj&�MD�(�/�0<�>��aY Fo����ֳy���<�D��8�94�1���*�F�+/@��
1�t�9���F�p$CnSNˡ��ZE3\�C�y�z��;=%�l��@,!����jA�Y�-Hpzj3�[KSjc�S:�;q1���u=3��ڐ|���Ƥ.Á���P�����ԅ�����Ԃ�F��6��4>p��u�S�?B#�pQ��[�Z�o���֑o�n�Rav�<�b�I�����[��5�����Cl�T�1	+7p��w7ݬ��bP4@6�
f��6��.Gh2��'� >�hTH�0i���.-T�A�l
7b��(r�
�9{K���۵�e�6�#^�D�������8O�����u�A�pc�� �>�����a�W'?��હ@*�lU�����V6���UX�
� �R�1Ԡu(J �R�1Ԡu(J �R���{�1�8 �[+ƅ���H�Q-�Na�AD�Q9�Na�A��u=�]Oa�S�M &�>�ZG�� ��$ť(���0F�-Q�M���-�� C��Ь o ��oBE��q;6���|�[��a��m�ϝ�N��i ���j�W����l�6�l �-<J �&���m."ゔ�RH9����H�&�!q��Ԗ��n1Fu>���`#�0��q8�O`G�Yj�Z�����e����}|�O��������f�3Ri5&�3Ro5&�3Ro5&�3Ro	�Ij�-@5%���=�����m�j�88� C����88� C����.$_Eċ踑}/��E�\H����q"�4-]����hZ���еv�ѡj�47��I�sjM#�RoړH�ԛ�6��;5&�ͩ7�mI"�Ԓ/�I"�Ԓ �Ũ!qj \Z��ÂD0��-CPC����v�����\Z��Wa�"�8$_E��/ ^�2�2��*��A���-��=�9퍇�c����%I�j� �-�D�)��V�[�7\�U�UnZ�$P����J�;�_���G��L!��1��QGTrG)TrsrZ��У�Z ��I�)2&@���� Rd
L�I�)2&@����*92c'Q2)V�+�Bc�RA��7'��c�"�Ě��)%!�$�I���2{��~1�h��+ঈ�GV����5�:�����P\S�ض�R�$��r�9ȖSsq۪ �sr��Gt	D#��m ��e*0�1\".k;���a#ТX��aH�@j�MmQ���GgB�0\Ğh5
&�$�s��+�J;�!��8LG���c��nT?�H����1�Q�9
�P��QH��qh52�%�Q�蛉����������h�Ev+�
���+�����=3EFZ�	G� �M|�f����۞jF�A`� ��I�.�m+W��l�m_��64P<�Q�C; �}<`�����X5?W� �U&FH-��Ă�
��p9�.�e�Q�S��
D�����-�9���Q5��\%MĶVZCqz��X�L����T��0|�-w?���w0H~46Z�)Y�57Z7-��?�ʚ��n���Vְ�i�A��Kw�ɲQ��!���ɉ�1���3z��1q\���U���x#�``� Ҹ����j�ư^M�^��<#q���l8��Zu�Aۈ�-��7��������C_�X�V��@q���W��YJk_!<.�6GSHCZ���ԟ:��*ԛH0"�:�/RM"�4�ʰ����	�ҭ"�Y����C�ER�H
�ɏ&����iGs�jO�О�<�d����+M��I=��)�ȏ=�#�=��~*�z�8Y�hwJN���|�6���!��Vy֦������+TT"�Y�n4�S�&T�$���qz��<�?/��t&�n�W͐���_6kŰ���*�[���
%���l �[zOBA��H9=	'� ��$����АrzOBA��H9=	%`�H�	��a6��,�{8�>Ie����Z�7��#�M :�=�ZG��H�o��E�;�G|�/�E�;io���j1�E>w �`�., 5$��jqFo���cRH�Q���������M��s��)����݃��1���ݰԑ�F:Ԩ"O:Ğ��@�?���r)Fo(�";�X%���C��_����x���ϝf(>mҋK���dhqm."�`��V�`��V�`��V�J)��E6�(�ҥ�T��J�SiR��)�ΰJ��:���X|���`q�$q�Ď88��8��GHドpX
|�O�`)�>u��ΰ���:�S�X
�O���>q?�'����8����|�~�O���>q �O�� |�~�@����{!�����8$^��a�"�8$^Ƈ���{OcBD0Б4-_�����#��A�DP|�8���`�"�8-APJ�J��ԯ��J��ԯ��!��c/c �����__�A���`[N{bs����{�-�rh7}\�{AA�pdKa�'=�O{b�+d��D�_�Z�-Ѓr�b@ĉ�R2�FFo�d�B�DP(�!@�(��)-pD��%�I�� Rd
L�I�)2&@���� Rd
L�I�)2&Trd�&N�drR�HRQ	I )	���NA�&*:�h�e�9H�DDe�!R��!C���Q1R�����\rhs��ƪ����W8C).5��Z¸5��h}4���-�H�y�j�D�מoG������k�A�[r\O��Z�E��e(���qA-Je�mj�	�tY�Z�Ja,����F�ӳZ�BM ��[�{�S5��JOm�� T�rn�S����B��Ę^��D&Ɋ�D䯂Yu�0�h�:����ph��ph��ph���4E����~vA��|�t�C���R&F��P�ր~��s��bCr�ԖmA�m�zv�W���H����E�/k��q��>��9M@a�&���l0@*�/Z�i[�̮����Ԑ'�TL�Tq��B��ÆE�:]��կm/��Jw�J�����<�"M1z�0 �-����y\~>W6E�&�U\�	�����i�-���x(��C#���Jbj���|��B���wq��0�k�tٌv�[U��+�Jb#Q����Z�I����Š�L&���gɥ F�,(��u�����E_��8~4�P�Az�;������ai���Z	�1�?������~:ڑ�c;S���5!`0��!���z��~8=
&��X/��H�rr{e�')�J!�σ���V'd�-��r\�L�HMDiz�74@��.7�f���SZ���V��6�N% �()�u@G{���PG<A�2PլV��� QZބ�C����F�O��"�����SL
�����kJ�0�����U�_���5�t:�i��̀��@:�N	����g�|F�}z�BA��H9=	`�H�iC��u�i�m#�M�s	���6��&�>��G0�H�4,�(�!O�D��8�5%(�ҰGQ�#��ciqQ�# �Tp"��Q�#e�ujyFZ�Q�FTgu�]��L�T�B�+�q4+�WΥ.��q�����J48�	Â�(|�8Ԕ��������Q��
v{�F��D��T�� &�4'���!q��u�^��H~�:����@;|��qj08m�7����Nn
T�[`�9��~�T?,��5���<.)O�S��n�\R�t��n�\mҋ��Qqfd\Y�fEř�qfd>ṁ�T����~�<�O�T���(~�J�R�����`|�,����`|�,�����~���������~���������~���������~������`~�G��*8~��Q����ΰ��H�`)��:�S�q#�u��ΰ8,C��P��GH�D��H�|�����~�2�>w8~���/ϝ��M��i�-6Ⅶ�P!PB��__�o� �r� �[[NNO{bx*��`�l�D�sM�`2��� �4�Z�&>�ܨ����:JK���Г%�p�U>M0���\����9N��$�D����"R�JQ�J9)G%(D�� Rd
L�I�)2&@���� Rd
L�I�)2&Trd�'N�ehR�������	Q(.��S��(52jU���е�S��$�RuH���]�lrZ���Ę�9'.:����Ю1.'���Kd�`f��H.�Y��S���KYS�7&!���D]jh�SuՄī��8p��'��	�ܝ̦����&Vi-yX��in��F	`�P�5'7!pN�3ڴ]�Y<�$���NBc�. RT�'�,�T�J�4 ��NDN<�)y�����$�����h�ƈ�h��ph��ph��ph�Ev+�
�쀴Wc�4^��4)N�@|k@>S_9���MIf�4�e�k;R;@��Y"�?nQ<Jj���ǩ�hչ�I�|MO��:x�Rn�CH��$aV�VZU�FH=��NX�G3ʗ#�h.(���$`�H���1��@��?�ê���,_6^�Q�uD`i��$�
��/W�W�M�L<�R�y��H(#t	�D����G�u���m���ҫMM+�iA���Zmw>�3���CJpɕ�""6벂i�:�M�_�-�Z�a0c���x��Z��iZ�L�M� �Qӵ&��6��/:gJ��`�q��01�M��@������[qjC�P�u7���apq�'����3i� ��4��*�I��e+�d���B�Y�&�~���y�k��m*��|���ټ%��4Q"D�Tዉ���+Z6�))�gSH��Ƹ"kzA��(�M�5�Os ��b%Oփ(#�DdƄ�j��\^�4��*G��ҼOC���<�#����|�S�-��q�.�XZW���Rc��L�a7S`&�P|��ϒ���v+�%c�uX :� V ��a֑�:�7��W��j�H�|���� �D����~8�/�G`"E�?5��t���`��26�_:���Y�	_:���m��)��`�pX%�
��)���\4,6��!�J�hm���QqJx>X*���͏Mf��5�W�ʥ~ܪ|�;oW�ZH��
���+�5��v�܆m
`M�L�-7���mZ}QԦ�!9ɴ+J1(Ґ;��u�ip���O.8������k<�q��ui���; �C���|�D?���Mp���h��h��h��i�D-�-7(����ܢ��Bҙp��\-)�Je�ҙp��\-,�K5B��P��T-,�K5B�͠ZY��T���(~�J�R����2��C����m�=5+C�m�=5+C�m�=5+C�m�=5+@��J-,JT����J-,JT�ҕ(��J-)R�M��iJ�Zm̋JT��ndZR��s"ҕ(�ۙ��E��ȴ�J-6�E���~�.�ˇ�2��nd?ṁ�T�ҕ(��<�ԭMJ��ԩ^��(��.-,�JQ�Ҕc�Y��5�;�Y��5�;���3�1�3� ��'=�[[NO{bx*��X���=�)�I����?L{�AGS���A'��H���%�j��IR��Z�C) 9&1hKa(��������I����hB�U��9B%(�� Rd
L�I�)2&@���� Rd
L�I�)2��&1:��+B��%�%�����<MTE:Жy������koCj`D"��h4��L��)_W�S�����l0_T%!�B��%�jk4ĉ�1�5?5�EF�i�Qeٵm\�D��Y�@��J";�������؜�ۈ���s���W	1�M\9)�ZN,�([r%�-����I���<yNji�CkkL$Wz��S���JO�'�i
�����$Vl/��!�SxMT�4�u�=RLй�cĘ������L��և��!&���O����O�$��O�$��O���Wb�; ���Ev=3Dq'��[C�nU>u2 �M���M���A�PЦc�۠m�C\,��\H��(�%�R�؉b�J��6�2xX��+����X�F�^�� �C���h�j�A��1$�)V�Zj�h/Tq����2� �Բu��C�4�րj3��po�GY���l������
#ર�B�*$Ď����kK.���ty�
 ����v�#�S[j�Ja{��>mD �׸эk\�15����R5��+��4���#�rE&�H>�"����&2�jj09(8��Lhc�G"ӭZ?7�'�"��J�D�!�V�x�X?�愁<.�;�Mʙ\W+��.'�A �u�ۀ:��Z�u��������x55������±��֩Ik�o1����B�P�����{xKI?�D����$�01���EGf���7�R�>|;�Cx���`T
�	���U0�D�]�x3A�䍀��Dp��D���p��(��lF� ����+«�A�V�R��@�P(��	��A�,�9���2A�FQ|���@D��"@R��#��"8j�Z���!J2Db���\E�J�����%(Ƥ�2Ԕ����RR�jK-IJ1�,�Je����pR��t��fy_�*��[C�m���p~�T��>vݡ�W�%~�@?5��\Y��Z��T�ەJ��T��h+���szm�驐zjd��~���\qY���?���ָ?5��s��ۗ��v1��β�A�cH�F:ے�u(��`��nq�68�T ����$�c�Ev��x�i^�w����6
�����ۮ��n�~SC�48SC�48SC�48SC�48608608608608; ��d��pܢ�A�r�8nQ� �\7+���@��h�m�͠Z5��iE�ZQif�8��+5Ê�p�\8��+5Ê�p�\8��+5Ê�p�\8��+5Ê�p�\8��&�C��P�kT8��&�C��P�kT8��&�C��P�kT8��&�C��P�kT�ۓ�ML��'��ry��&�C��p�\?�ƴC�P�kT8�Ҏ+4�����k8�����`pk��A���'=�9��lO{bp
{��S�Z`��Ƙ&6_P?rh>s\|����U�Z�s�'K$�k��6�qqȈ�䄨�N�I�6C&�D�(�%d2Z9�p	�I����r"�DQ�^@�(���R�
R�JP)J)@�(���R�
R�JP)J���Q2���B�hR��$e$�%N���[�D�xNhV���(��ʔB$s`4`��(�WX5����J�5�#�U1���)�j���v�vl��N�w&��\V;�)��kj�1O�喚�N(�js'�)��a�w4򰜹�RD9"y�HIuiY�Z�p��@����]N5*_�H�F��n�Ddy4~�Spq,M�0�]�8���#��	m�5*QR�Ij�d�J#Aǁ]R�$��D�i	r0.xr<u�W ��`�O`�O`�O`�O`�O`�`�`�`pO@Z4"���B!hЉ��BL͍
��?6 )��87,|�dA�r��6뀋A�,:������J���hn*`���4(�!eb�u :�<Z©Ma	�b4��@:�TWjJ#�:E<j�N�A���.@񚤭�6ܛ��*Ԛ�'�6�`��V��֋� |^5Dm"{��OzG���ADn�R%A�DI�4��n�;�m�Erj��`eV*�����u���:�����|ڋխ��mi^'G��>�[�Hb}]sG\n��~접6-Lv�-<�8~9�@�#:���8�9֣7��n�h:�p��u�������Ai��jo�hxo�q�Z��d���@�?��c~�GP��Lw���c�#�i���w��W�3�Z���o���CېG�j�� 9'��ø���Ш��^B�*�"O&�4Q��R��Hk;�/^�16u��M �-dƼ�a��hT��#��#�8du� V�ecz�/���� ���^�(z����CАj��[�M"��4�A�Ip��}���m� �x ,� |����Tp#x1�Z�-N� �S�2E+iH�m)-I�q�,��B��аJ.6�E�)�q�J.)Oƶ��f�>5��5A�>Y��m��+���|ۙ�s!��(��\�ەA���_�*��[@~�T��v��f�_��=52Ѳ�0�M͈+󲧦lT8�*d�?71������
hp��湌�ζ�-)�aq����T����
"�	���LyR&�D�HM��QX?I�����#�85����^sZ9��l�wb��WG���>SG�Z�Jx�S0~SG�4~SG�c�c�c�c�c�c�b��؀�l@~6 ?����������������2!�L�q6*M��b��بq6*TȌsb:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:���r��ܠ?�(���r��ܠ?�(�dC��P�lT?���C����D?�(��Z��Z��Y�L����72���h:�ǌu1�Ld�S1��\�1l`[ �s��؞����'��=���i�cL/�6]�|���)���<ط�[������SJ�&!�� �$O9	�R�G![�I�99�R\�M����.�%�D�ФšJ9!G"(D���Q
"�HP)J)@�(���R�
R�JP)J)@�(���R�
R��(������Q�H>J���O�bA�[X7���RGjd��Q,�\�5����`��٤PS$D���]`�X$�sJUM��L �mK��J�F%��nP�4�mV��n�	�>(��k���}:)E��Z:L�y�N@
"@�	.1�K����b���SS_8
�fȐ������|F�rt��9&<��Ϗ�@»�Ũ5�b{Y,Zr��LD��&��I�eJ"ǉ\PD��c�Ev��IsĄ��Bcp�p��	Lp��	Lp��	Lp�~��lq	0q	1�����B'�O@8	08	1��EuϜ���M����v叝�ciR�Q��T���XC�Z��@hR��˟;r�hR�8���p�X�(�@X��/�=��y�Q�G�A�Kt'�]��A� y-���r�mSr˼��v,�Z��ɬ�>�.��&�4é�A�p��V��n���So�mzBm�Ifh����mWyB`�e=.�&�:�k;��s���mE��^w#B�ѥ,������V�Jd�͗��4�K4<W�R�"�o)a��I�5�0�q+o���F��p�!�����u��7���V(�#xJX,�x�F#�����@��h9zjՠ�Jy�����Kh�͠~6��,��hC�Q�,��o�E�����Z�������J@�[^,I����UhBZ���꫐AA��>Q֊dӼ��l�[ѳKղ���w��X�B�hV��m��$v�ꌊ8���9���IN#�$>c���AN�+ª���#V4�j��x�/I�W�5����<T�!OB�`u�2H�-N6�����<ԜJ�e���Ĺ�q.|�K��UͥJ�\Y��3Â���۴�5A��P|�T��k�9�s�5�۔A�r�?nQ�� ��D�(���~ܢ۔C�]�6*�iC�ZQiL��=3b�iL�_�*��[@~kh�j��r�驐�N�h��צW`�h\?�f��YهY�u�#��?����8����?��[s:���l��x�WD?��s-�Ў���`����Px��2ZɅrk���P���"n�&�_6���������f2���R�M��=(�"��(��2���f�h������������������b��؀�l@~6 ?1���1���1���1����������!���+����#��ì�:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:͓��:�莲�#����+�:��:��n&�q6Z������vcq;0�;"jf��Lع���fÇY���l8u�9����� ���=��lOOi�cL`��}A����9���:<YI��M�Zq�N~!��JM
9	�
"@
L�Iq�:���A	��)*Q���!��R�	�a:�V�x�E��R�
R��ʎL�JP�J)B%(D����"R�JP�J)B%(D����
R��(���Re��n��J������=�F��.K3
"���iֳ;�f�5�H1��ܩV������Y,���qH��q�'?���%��i\M\�p��WC�5�|�GR'DDMi�ٯS֤��iH�p)*1ɌHV�"�At`�&���e��"mT��h��4�u؍���3��d�eHH&T�܍Z���<kH�$��qв�l?^\�sBrФ��;�%�Σ����͉U����Wh^*"]R�E{q	Lp��	Lp��	Lp�~��l~���zLЈZ4"zd���lq��>s��dhnc�s��~������6�m�3sQ�w�Ĺ�W#�N$�dpSB�A6�PK��\�V*
�=Xu�z0�Bԛ�1�9��ZX���X���wyAzPZ�5:�`���'�AXD�6��`�H�U�Т�0&�rm����Q�/��-�'R�|����$>i�1M�/�A CjcSJ��i3h1�׃-���6�_�A���zf���:5Q�!������F�Ö���`�X8>I�~ԗ��iw����q�
0�Z�����c�P�?
+��B8� ��Ha����phBm��4�8|/jO�����
;q7� c���-���b�0�|���m#����m��|���
J�I��*fԀ,�&�� ��~/p���bԬ$]< �~CFI�8I�S_����m�dHZV��U(~�4SD�����8�A��O.~ ��Q֮,�v��u���4�pu ��:��m#���>�TN����n�:�TH�-Q5'椑@hX"����,���xY���lQ���r�\6|�ƀ��D�,ۖ+�5_���M��h���h���h���h���h�ì1��⺡����'�:�Ha$sB�8S4
f��\8��ff��O�xpW�Ƅp���hjd�ML��S+�b����L�jf��h�2����1����W����@�n ��L.e��6��s���694�R�潁"hd��1�hi���ե'��M�Xm2�,�n.#���Z�n@:����z;S�D(|"��y��I�je{q;[���J��W�����įn%{q4 �M7B�Ѓq4 �M7BY�u�'Y�u�'Y�u�'Y�u�'Y�u�'Y=�Y=�Y=�Y=�Y=�Y=�YهYهYهYهYهYهYهYٍįn%{q+ۉ^�J��W�������n'kq;[���N��v�������n'kq;[���N��v������Ѓq4 �M7BL�je{S;Z��c�L�mkh;Lc�#��;"1��A��h+�mt��������ll9���ୀV����|�j���kw���#�R���	o���rsC��!�o92�U�yɒ2)@�$M���G'"Q��n$�5��^�G"(�E��
R��ʎNb�N`����"R�JP�J)B%(D����"R�JP�J)B%(����
L��b����"T��;7&Z��Y+Hca"rUq8RL�аYQ�į�@%abD.q�S>���u2�l��o\M�jRZ����	�!��H#�^�&��M��|y��H�ܷ�өJۤӹeȬb2k�!����C�2���Q6�%�$���jVݯhV�Z�:p��<�I��;[�"f��md:nT` H,�!rkB��S�D�"�]��'�����"rWZA�ɸ�Lpi�~ܣ�M��lGu�۔�rv��q�~�~�����Xc���tC�]�@~4 ?1����I����	�Ev�h�ܰpnX���M�����ҳ���h;Z��X"W��`y|0<�2R���D#Hm-�e���\QBQE�$\5���I���cA�Ty*%M�F#O�]�)�E��@1hj8@�A==�b2?,��xT�(�e*a�Rs1ۑ�i| ���Tp+prri���Ǔ�K0�p95�c�˾
�h�rh	���U�zu���
i�x���FV7�;x֔>�I"'��LH��x�8G��?@�����;q	�Leq��X�yژ�9:�:�u��������c����x�m���hW7&���x�Ɛr+����
���&u8A��k��֊8�y�;�r-<"��"�ۈ~�#p1��`�J%ͩ��67�a7Y��S��� �M�V�R&��(Wm����Xۋg�=�Zב����ҀKC�^�/M�"4��DyV�B�]c-�=�;�k��ZH��5r`uD��:����M�`e��ҽ���<ԍ�b��q q[K�Ԗ�a�q��&��,���,���3�b�]P~vT���=52ML��l`�lc�;^�����h��h���������dA
���$��A���:�L��Q�蚙]+S+�:��r�����'��gP6c��9^����=�"O<'�m�M�Љ�	^p�G'Π�G'Π��gPJ+��y�O���7���Bh:�G�a�Ysp&%�+N�o�y���;�p��e1�����	-�+*��D-+	 wz�������A�pv\8��ML$����O������)���)���)�a�a�a�a�a�a�a�a�����O������)���)���)���)�a�����)�WD�NȎ��&�vDu��7�#������7BL��q4 ���7BL��q4 ���7����įje{q+ڙ^�J��W�����įje{q+ڙ^�J��W�2�L��S4"jet�]�WA����1���mtA]�W@�;"1��b���v<�
�[A]+h+�sv����o��Ϸgې*��+l?r��H��͛��oJ&$mXi8��x���>
J�D$e$%+�B��*�B��+�B��+�B��&(�&(�$r�rrr�!Hb)�!�$2d�L�ɗ��y�ל�y�Ly�Ly�Ly�Ly�Ly�Ly�Ly�L���"R�JP�J)B%(D���R�rB�I���Iˇ$�O�ʹD�1Ίf��j<ۓ�$�D�t� 5b����Gx�(��a#Y���ZשJ��bke K>7�m򝠩%#oe2k�`$vR���CA8�PK+6Rh�I��z`ֆ�B\��Ed�S-�X3xY{V�͇G4�����<�j��n���Z�
e �]bF�P��`攋r�;�֭�<��v'-��j	b��.�V�o�af9+�$��
w����DI^
'�^���C����p)1����c��q;
����=+h�!y%��L������Ѐph�x�W�Ex�W�Gk�nX��q��v���Ksq����靡Ղ�b��yJx&�<�M��&�Y��M�,��%�Co|�w0j��3T���'��%J)1��i�.j#8+�A�n�Q�ө �N�����":��O!��Tv�dXښ�����		�D���k��p�J��VI��.N~J�!,A�и�|և��@���V$��'�U&�:e~�Z)��ڜx�ލ-k[���࣫G/L�1��[��LeCW�;q�3\���-gP��Z
Ј~�%=4��8�BS�x�EcΑH[v�hlY��D�Q,.��|�������m�ȴ�%=7���ա��_(����Cm��7�E�m"D�i%�US&��U�:ےDBD�hV��R���hx��Bѹn
c�du��H�R�]�6����i���- (��l�&�,T�h3hb�mh�y-"48X'� MI�q�q.�Xq R�6�e�@uf�:۠�,�Σ,�A�8,����s�RSE�4>S_9�-���Įì�:�������������ğI��%�������Ё�OD?���C@�1���B���uĢu�MDGW�2�Хr��DH��F05h�:�Q�R^R��>a�#����
J��*��x"h�
RQ��A5Ğ1"�
�>��f0]+h!n�M�.��K��ӁbQ�]*0DqXLJ�4�R��F#�<�]�'�+�ID���<� wh���	�r��h�B&7��/�m�/n&7����D��"cp1���Ln&7����D��"cp1������@�����@I��$��a��@���@��@�Π�P6uj86uj86uj86uj86uj86uj86uj86uj86uj86uj86uj86uj86�Ln&6���I��$��ch	1���Ln&7 j&�cp	0
Ocp	0
Ob���+���+���+�A�����(�%J8IR�T�
��Nv��ӝ�o��p	�|��tM���Y���]�M.M�IЉJ�Q �&<�+�B��+�B��+�B��+�B��+�B��&<�&<�&<�&<�&<�&<�&<�&JP�J)B%(D����"R��&<�&<�&<�&<�&<�&<�&<�&JP�J)B%(D����"R�JP�J)G$�Iˀ���99D�ǈ�YIS��@�|)	�x5ɼ1Hau��M|KT�W�<JǕ��&���Y�,����Y4�:'RO���bH���Ӎ�e���0j""R��v�b�+�I5�@��1x��LFA�Ԥ��\��O;��C��Ҳ�̠��#������st'�J�Ta9�ܩ���ԬH�S�
C�ad�Nn�$�u0I�S+'��O�#���q�wA�;jm�Lr�n����L���»����ܢ�#��q�5�d?R�|�㐴�rm-�dZ'����")(%!�&1>c���=��=��=��>!��-�-��� �M���M�qM��MJ�����@�`t���� �؀~O�V�k[RXE��hH0F�D�������$�̡<0����Dd�eҢY#A�!�F94��ئ�i�Lm�;����l1h�B߁��?��z5�*5<��GtkhS:�1�����Dg�T�`�X]N�<
�B��V/��S�B�p:A��-����R����@��F��c�'��qH/�Mc�����������p������a�&�C���?��MFW?ژIL�&�M�x�Y�_ˈإxn�����HU����+�����u�1���o���xa�Ԛ���j�F�Q���_����Z*Љ�@`�Y�����Y�D��L?o��]	�R׻�$�+B���mT�sh�؉N�'8
�+6�
��ש� �]ڨA�tG�ҿU.pu�ѧR���S|� 
2���	�a7�Rړn��6뀋4�6p!��[��k���?na��͐�M|���;1_����������jf�S'��	 u���H�$j�I��6c��8J�BV�Dc�50�A�h%gP6c���mu�85+���q6N����v�)*�u�79	�QA>��kB�h_)��淶�W��E<BH�F��ҎI�a
�Lb�8�h{x���h��L��$Ä2p������rZW����N��K��%K��4��L 9+45r�ʹ4��u|Ln�I�j9
�W���4^r����G!^q���H7���p! �H7����Rb�Rb�Rb�Rb�Rb�Rb�Rc�B`D�����!^r
"`D�(��Q �&DL��0
"`D�(��Q �&DL��0
"`D�(��Q �&DL��0
"`D�(��Q �&DL��0
"`D�(��8].��AG����Q��(�tp� P� (I$�
D	"��BH��$O85���A���Py��<��pj Pj�(5p�
\�����s��|�"P�&^F��$�czũe	-p8�P䞩�+��P�J�Q �&DL���9
�9
�9
�9
�9	�9	�9	�9	�9	�9	�9	�9	��"R�JP�J)B%(D����"R�JP�J)B%(D���2d�L�ɒ2C&Hd��!�$2d�L����n�ML��q&�A.��Z�l�rn[���̐�PnJ�Q��Jл�Ef��X7M����p]��B}I/呫�ZjN_�oVKo$���iͯS��@�p��^��5?�
�"j��kH�Σkx󄖏b�$�'H��"�;��@\��"(Y�VH�;�"�(=�ڡ����$ (L��ԩ�M�$�l7!%#�N�I-�B䍗�r�H��iD���h0[
b�wQ�%��̼�d����$�h;9��E� ��m�"`�D��m&�#��Q-��!��{1����	)�N`����Dì���!0�ژ^c�Xc��8J?��8��8���]��^-�����������?�����V���t��� e_��.)P�m�gzf�~۠��k�j&���U]��2�p���i���56��b�@D�4#^����om5D��p^7��R�LҤY4�΂m�dy��C��,_,��|Kw��d��v8���%r�:�#:�	h��@H	A�������B8ـٺc�"�� a�?��MFQۈ�o������|����[���� ���3�hx����B4+�c��u��-� ���w�$���U��&�n!�.(�3i��`�-s�hyΡ�zb1��Z�p1�������4-u~J�Jti�ԲHH �aЪ@l>5��M��@�P��q� �`��p�B��Є�4��H�d�8�٭$R�\�6����e�y�)�v���G�4*b�m��l n*S����b��RX_'������h5#[c\\nb�s��~���5�"��-��^-��]���#�>u�'Y=�0Jc�05�05q�n ����)�����mL1�L:�HE%J91rЛ:��D��m$@P�ǜ�	���֊g׈�����:�HI�Q:󓣈68��Q9���� ]SHh.�4Z�W�w�	<��JH�ZЄ��'��B�ڴ�Z�Bb$a5r0��NJ)
Z�Iˀ���y�ա9s����K�1WO,ɨ+TMөjD��)Im5�9���r�Pp�G%�:��c$(D��&0"L`D���1�c$�<�$r�9I����RA�) �y�L��BuhN���Q2J&G%(�!��C!0�Ba��	�2d&�L!��C!0�Ba��	�2d&�L!��C!0�Ba��	�2d&�L!��1�"��R�CHb)E���"`D.��]��!vB����"`D.��]��!vB����"`D.��]��!vB�y��p�'�.���l�Zb��S P6��F�Ф2�5_˿��_%D�j!�69ւ*Й��9
1G����Q��DLy�P�J)B%(D����"R�JP�J)B%(D����"R�JW��ǜ�ǜ�ǜ�ǜ�ǜ�ǜ�ǜ��2C&Hd��!�$2d�L�ɒ2C&Hd��!�$2d�L���Q:C%�%�A5�5D�F���S%�r����QǒI۽��b[Y���D�w�Il"�*F$�+V����;'�ƠH�L��S�??�F�����`�ԋ"q��`�kN7�¥�Lb)�ZmS%y�H.�S���Sv��`�^:t;,��T�8�@�4�F�MTth�'�e��L z����i�������6�<��F��j)�J�M��`��@w>;�ަ���ԥ$'[
��y�R~|+���;1��M���F�;=�	�������"hQ�	Z�])�h<!"V�ش&��F[�,�5c�M�I�Q�H52r��KD�
Lm)�Bcq[��u��X^?��I��>��>-��>-��>ua��-#��.*3n�Zq%���ep!h쀸h`�?�I�`j9(��n��fy���T@��6����SCxY6�Ԑ��5�\�1����驭X�Z�������t	���P����+�K�b�$Ăj��~�z���7�Nf�^$�6ҵz&�QP�۵E�Ykh'�E����R*u�d���**[~0NN�#���9n��@�V��- ����|�;q��*��y���j;qF8YGn G8��xm��|�K�&�n+��SH�-ʕ��:�+@�~?�1q�j9��^s�h�����ͤ�1���~	��;�n�p�ޅp
���/�śn6�NZ����ͽ�E���tpY�+��m�b- �q	�ʴ.�m)�uX޾t�ZܩڧB���A�x�Ē""LNT�����ǚ�T�G�40��lj%����M�iJ�)��\m����qh�Ǧ����71h��צv�x�W���O����O`�O`�@���������L/:�S�E:�L:�L1�L1�L1�L1�V���)�"�G&@��<��D2Z"Q9����n�p& 9&"F����$"�1��Z�QI�š-��kA.u���j��j�DMA"LT�!uA�OjbX��H3S)V��B�i=�&MG&�����+I�	2�	1���IB.�+1�M��)�R�亴ku�Q(�'�`w�]A�Q&-*�X%�Mɷ+��O��Z�a2�!V���S\u�-	lF��t�N���:C'Hd��!��2t�N���:C'Hd��%��m�K�	ա:J&ID�(�%#��rR�JQ�J9)G%(�����rR�JQ�J9)G%(�����rR�JQ�J9)G%(�����rB�JQ�
9)G$(�����rB�JQ�
9)G$(���2b)���C!0�"��L!��2b)���C!0�"��L!��C!0�Ba��	��Q����։�K�I�+��������L���PJ��o9
9)^r
"AG�Q��p� (�����J)B%(D����"R�JP�J)B%(D����"R�JP�J)B%(D����"R�JP�J9%�$����\rK�Iq�.9%�$����\rK�Iq�.�&�9&���XcXc�1��:�����n��i��!�ݤ�"�D�⚑b����	 ��_r�mjk?m��av�Q���o��9�@�cn���Nw�K����L:��b!'��o�c�����t&�����Mi14�	ڭ�����)[����59�K�*8��$k���yHF�(_���g�,��nWt�M��StM�i5�5��m�x�9��9$"j���
"�|�i�F�J�J5D�;�k��Fl'W5�),c��)�"u�7sB�b����ZC&��OF��eik%��<��O8� ).'Trd�&N�e����jd)���x���x�������y�O@q5���E�f��.�D�?Y��!�A<`~�֥�����`RkZm73�h]<�v���e����@��b$Vz��V�#Wz�LRI=F߁#�O�H��9R�	#VC��3w�4_��u�<�Շ� `u��&�fR�7vT�+�
R��E0F�j��v��W7n+���Y-n)�RoH ��eo�r��jo�q����OLr�j8��!��Z0�I�[��|��TD4�Ÿ�G"�A\nT���u/��Z?<U���DC4)�ev���i	N��pm�*֑X󺗍��uV�ѷH�[�PE&�ji���x6���G^$�#bD�47TK��5+N��L�P8)D����P��-Q��=�4,�Kn6�+��i0Hj<|�?6�7�Q�3���G���ǚ�hJЉPf�5�?$"��xZX4���vJ���+��-70�M���צ��F��h�f��h�}���Lj`�Sژ^���D��Ba�B@�! �
Ln&JP)J)@�ʎL��ʎL��+p!Tr�G)@�������MT��x�`P���T�	�(�$�wQ޾&�u��e6+F�)1�QI�KAZM@�о+Q�Y�V\�+��F�%f��4aI``NS&$���Xd��S��e�R}_�ք�ui�rК�ZN8�;��)�?��β��YN��$��M�Jw�6�&�݊m��xHu�� ��f�9=j�tF�jQ��Y5��Dk1�K���S�j��M`96�&����|o�m�M�	��-�B[��-	lZش%�hKbЗZ��u�L�	��2�)1hRbФ�i:�'U�괝V���uZN�I�i:�'U�괝V���uZN�I�i:�'U�괝V���uZN�I�i:�'U�괝V���uZN�I��2�&_���|/�e�L�	��2�&_���|/�e�L�	��2�&_���|/�e�L�	��I�B��&-
LoJ&"�-���K�)yɋ����B��+SL`m�o8�9!G$+�B`D�D�D�D��B`D�!�$2d�L�ɒ2C&Hd��!�$2d�L�ɒ2C&Hd��!�$2d�L�ɒ2C&Hd��!���\rK�I���k$����.J�D�(k%d���M���P��)�%�JlnfJl%XM�Iv��W�����f��<��z�6��\�Y��֌	�ە�i0��wmF���Hf���҄hdidt��׻���q��X��SkL���?))[�r��*b���y�PIޮa��;���� j�b�ڟ�-'7�7ZͯR����()�$Ųi��|��`F��S�:���"4���R�᛫���VbJca��� �S~|5��Ʀ�A�����!#���Ʀ�W:.i
`�5�hi�	a�%���_!�a[@9Mr����ib��%��kd�#U�3J��5���<�������n�h)Z�J��S��:�S��1�V�R�HH����q!0!Z��`�O8����k�'�1͸��e��1�p<^#cr�0"~G й��E��������\�Ѣf��z��$����ޤe����"($Y)&7Vʚ�u��m��)���ݾ��ή7:�.c�H�������1��O�W+��f�	�#B���Q�����P\��r_�(r2P���RKSY�W^*����/���:�h���:���X�:�t������3����Ʒ[n�V�JIZ��WV�"E 9^?ښ�r-�w�9��9�4@��E��X��7�&mH
��p1����F8\W�Ch1�;q:��H��G�M�@�ZC&5^��tpq;�Gr���O�IA! ��F8�	��ly��Ցtj�y5��4��}*��iZ8])��  ��l�Y������ܾ�jds���;Ls��+ڙ^���įJ����m��P�u���n+p![�
�
Lm&D�D�D�7j R]�'Hd��y�ל�y��).�\"K�Ir:J%�Z����BjV�5x��!��<�rb�aZ�mk�$�N���[�N�����x�:�IT��7�T	E�GQeq(ă�Ă���b1	>E'��ئ-5��$
�׃Q���d�4М�j\S2�&�q)�C����%�I�W<F�r�Y��0rr&�ܧ7��n�H�ȗ�'�a���:*R��)
Ȗh0;F/�ȁ�Љ���N�ed�6<F�`֭)уZ��Fjҝ5��&�V�o��ɷ�Հ�ڴ��i:�%��L�	�>	��1Ф�`֌&уZ0�Fh�m5�	�`֌&уZ0�Fh�m5�	�`֌&уZ0�Fh�m5�	�`֌&уZ0�Fh�m5�	�rl�&��prl�&��ui-��uZKb��V�ح'U��+I�i-��uZKb��V�ح'U��+I�i-��uZKb��6&�,UK���c�8!"�㒜~4[�Ju���NA�KA�MT�&�!��<�$ �$@R'���D���.J&�d��!��2t�N���:C'Hd��!��2t�N���:C'G$����\rK�Iq�.9%�CY(k%XJ�CV��PՄ��hS�
u�N�)օ:ЧZ�B�ZVAhV@�V�J׉Y�j�"KA�'R"%�@��j�O4��V!�@g�K΂����OmNɠ��$󢑠H�jk\�E*IDvS����^&Z�l���N�҄�S����Ȍ��l��ko&�ͼk�&��ܮ|�tN���6�8���o�e"�ݡ�>����Hωi$i94@LoZ�y�0�䭫e1�S�^rY��<0��f�b;�x����V��V�M�ꝭj��'A��?͆	�:��)XNvY�^�gq�"�0��V&9�E2��hDnt)����[�M�D�;��5h_�K�г�`R����+^r̆V�
q�ZC)��Sakyɬyɵ�è�:���1���n$ɌN�V�N\cmĤ�~;
p�����cq;�+ǓZMi�N�Ҹ5�M;,[S�hm�D�p��Q�U.�D�/D�(�d�u1�)���ů��
~�l���	$�M��I~|@D@�#S����@���$A���c�[-�J��\G���4Г`��u���Yl��p�؞���gR��/W�5}m�&��n$~1"mMN 6�'2L�/IC�~��8x,j�#�zb38���h8À��U�T
���r--!��r-<U���"��/����Z�����p�ژ:�qV�.[Su+ ��r��Z��é��1��JM�c$R���c�q��1�H|����ژ��^> ��Fm-��5��WQ���+�&�{n�>2�y�����:��eM���,
����j<Mt	��ԑ���t=@߅=�	^�"y��9r�M���Hu��8I��S9�0�������m��O����O�Az�"��*�B��*�R��ʎL�����).%�%��X��Pyɬ��B]hK�I��X9&�"M`���Z��ڴ��Жy�K8�'Z�8�W	er���(�!���1Uƫ����5\�4ц��%�囬҉XN2ܓ�)�G�gtO�j��'�X�D�e�4��_��MY�����»a&"vmͩ\$���,3Hנ�,�I�K����L�	jw8�5*uPI���MXY�
h?��n[T.04�ݔ�J����b8l�j��$�+�E:�'��&�2݋C�
�Kef?�w�Y���Vc��x��)х4#Z0���kF�x�h��S�F������<	��5�m�S��w�N�)��;������S��w�N�)��;������S��w�N�)��;������S��w�N�)��;������5�F�����#[�kx�o��5�F�����#[�kx�o��Mc��xX�&��<	��5�m�Mc��xX�&�d���rTa-R0��Q6'@���B�D(�%��m�5D�%�?Ƀ�C���2�9II �1��t�M�F�:J'Hd�(�!���t�N���:J'Hd�	D���(�!��%����M����6J��(k|d��V�h�V�h�V�h�V-
�+Ju�YiN�+ �)օd�d�dHB��
�ܚ�O%�ɋ�N'g��@�i25S�׍�K�������
-k���� ��j��w�p$��G����bF���� |b*.�`ڝ��7X��čC΃I��Mo�[�|�b�5-��p5���TOS�����Do�ǒ�=5$P���m���&��ZZx�`��Ut�� R-�*.�s# ?{Lv>*mI�F�`M4��[S�p:A��k���"<YX�)�C����T�i�͵6���4�ӿ#WF���\��i�6�+�g�����V��Zi�Ʒ��ǜ�%��K�,|�Z�Z�%XC)��5�� �� ���.�	v�N��]��R�q	%zd%É	Sh!nM�Y�=ԛ����*56S�̩
��e7x�Ű�~T����{=ҙTx�F.T� �L�̠L��;'�L�
I	(&5I��@�^҅���^jX�Mj���QۓkSS)�Ad?�G����c6�J`���GT�C��O+�-P�f&u����#�jwW�0��`hl2<`�l%�ț-� I��B@r�W��q�&�n-�"�q��BRA\5��ҒE�;���uq�f�	��sB��KR���j��"mMEr��'��"xR!7�s���W_�� �5D�_7k�8%U�"��o���V\(���Cm����8|�ŧ���H�zo��&�3��H@�jM)���h�l�+�M��O%\�{�
e��fTm�j2��?��*��rj&��jG�����s@m.�*T���o�:��c���9ٰ��j9<2�J���@5p	1G�u�XJu��8��R�
R������Ru�'Hd���D���� �M��%6���6�&�V>�|��h�V#7���)���%�|���
Ґ&�\�+FW<N�i��mj���&�/
k�f+��1U�{��W�H̷�5�X4R@ԉx��e�dӉ[��j��n���b4�Ml+TD2a\蹤)�uF6�A�hW����b� bvnZсu���B@�e�BJ�)��mfƾRk҉�$�\�X�e4ry��H.�ho���\�)Xj<�;��;��v/�,V��4��i��Lu�n�f����Y��+"x��x��<Jh<JȞ%4%dO�&i��7	Z�4�e;���YN�+1�S���u���e;���YN�+1�S���u���e;���YN�+1�S���u���e;���YN�+1�S���u���e;���YN�+1�S���u���e;���YN�)���%4�[Ħ��kx���o�'�5��'�5��'�5��'�5����SA�5��j�a5r���Ж��.9'G$��Z��u�Nc������xKT�%�F�V�ش%�ZKbЖ�i-�B[��>	�rm�M��o�l�|`�ڴkFjҝ5�Jt`֭)уX9Z�)��ׁNV�
pr��V�W���11�i�Lx�h�&�������b�7���,�%��������SA w��H6�'��պ�W5M���q��a�Q��\L_ɏY�4��1%n�ה�5�,����à%"I�٬����dGA!E���IDם�*D�5�$�!�z�O)���
 jFꑭj��E����I9/�R�2s��b[PhD&�D�'��,�^��4x�ڑ	��c`5�k7�P~��.��bw�x�d �$�g��5����X��Ƨ hհ'&+�G��׶��bM8�۾p�9e�֐>I��հl_�MG�"�:��R�?�NJ�hf�ҹ BGm�H)[[��oZD�o�0��u�HEօ6�a����d#UÑ��Y�Z9+B#XDk�j8Պ96��He(�R�DٌY���N�d�$���"��<��~b4��>~�Uh�!T����Ud���s���òce�ש���)�yU�t)E2`���kU�P��k�r�|�,�������ZW"n&��Wl�e���%�!����MkL>q(���|����pzbEBm�e�����R��U@��Ou^q��:ê�R�x+C����CJ�������|�����@)��^�~,E����7�c�"0�hiGi�[g�^�ڐ6���R&�K�K�����8�L*c�"0)��U��~�|=38� ��e
W��i��I�R���FjS���y<�Dnn���SS)N���Q0{nS*�C����-���Ц�>�[�B��$H&�R�z� X��2ZTJY�ք����%��B�8�B8�J�[�]Q�Tc҄IӨ���Q.�%�d��N�Iv�K����%o�m�5a(��"N\�1V�{p&4�h����;��ǉ����bc���	��6��O�B�mM�7Z��-jUq�c��ЬMW���YAxVhiLR���[p���-(����3CHY<ܛPW�/�e�C�$�8�@.��&�o��D�BF�q���^7��d������&�ܶ�	HRE�bEd���DOw�q�M�؈��5k�[TF�Y��5�jLۖNZ��'����]�XZ&��i�m+�I
�pM�Z��6�^�^j���Y���q޼;ׅ���^kýxY���f�1 �,Նڱ���T���;��z�W���\b�5q��,��*L�_i3|i��U�1WƚL�_i3|i��U�1WƚL�_i3|i��U�1Wƛ����Z�4�xV�M,^�K�k����Z�4�xV�M,^�K�k����Z�4�xV�M,^�K�k����Z�4�xV�M,^�K�k���L��YY�M��'���j��M`8Հ��96M��om�M�I�x�X�&��Mc��ǁ5�ljǁ65c����M��X�&�Ƭx`�V<	�q��<
��N�+1�S�
�����;����N�+1�S�
�����f?�7	f�,�%���p�o���Y��7	f�,�%���p�o��&b��{xY���q9�� �+��aqA9)���"Yho���x5�5��S�����Im�A<�(D�8MI:<�<���k�HK7,�%��
KA9�X�W���̄�~45�jGxe#^n�1���)����,����yA������&�p�M��j�6MBE���k���ؽ˩�'�e ���l�J ��4�H~6�>���'/��7�I�~�v��Mc�!QH$F�Z�Τa8j"_I� 9Y8LI��z�Rd�I�ڔύ4���]Lta����_nF��D��P4���S;8����m�mc���8�0���;��w`9�iY���҂Ь�Ь��!��C�%6ɰ�.���.�zd��a��8���[�����	�%!-�(k��&<�0㘪9�B��� �T��<���t��v�I�R(-� 1���n�6��ղA'��F%D�#Px����J�n��Cυa�|ܽN��q6	�2��FVz�B�T�A�[�/'��A��"�@hi
��dw�uC	ڣg�稅%�,������&��5"hD5'$I�d����+��m�n�n[tb�f�n[tcn�|)R+E*Eh�H�M����VRS�q��C��?��:���׎��H�RRE�!��'�`�%o�r�S)A׏�x�р�����o:�X�H�*�`By���?,���r֑��p���cC--0 l&�����bpгOzeu��Z�1T�����Hl��V�U�d�j��OK*C�cr�y�c�2�M�[xߖ�ÀQW�6��d�D���V�B+��%�$��N�Iu��c�����Mc�kx��1V�)���Vc���Y��11�YA�YA�Y\�,��mj�m�SJ�+%Q��탩�0q��IR-jWSj��:U�J��A�5*qQ:��UƓγ��ݎ֬k�&��RW���&�*��]"Yh;آ+�����k�:W+�cj1�yM��&�����om˂�1
Z��Ro���V����V��$�B�`��%�����	<�jj�HG�#�Dj�i�+v��h?)��V�h��Zy\jA b���HY��5q޼;��z�Ԃ��^�W��R
��Y\�5U�mDm��V+���a��5U�z��V��UXw�Uaޮ;�Ś��Wj�\Y���qf�;�Ś��Wj�\Y���qf�;�Ś��Wj�\Y���qf�1 �4�xbAxib�Ă����᥋���*����,�|b��,_���K�$��/H/,^�^X�1 �4�xbAxib�Ă����᥉2�	2�	2�	2���5�Ʒ�����4�4�4�[�kx�hS�
uiN�)�#[�kx���o���SA�5���u���e;���YN�+1�Vc��p�n�&����	��11�i��Lp�n�&����	��11�ibL�^�3Uxw��U�ޓ5W�zL�^�3Uxw��U�ޓ5]E���S6��ޮ)^ܒ"'0i�a-�ALjD�5 �,�^�)VPk�vp\F����+zAo�䶼�	�J5w��IH� j~i@�٥4)HYN:� ��U#�H��NS�$0�����琛j6�6�q͡؁0H�޴��8����䍓<Ҙ�.~�t��q05�Z1�j��Vh°�5J�t7-�C��T$�i��7{(X��ܓ��>��F��:�,�&��۸ImxIЧ�����D(.$�ZMɤ��Q����5_��oU4���^����BRNő�ssa8�؞�+��M���*c��)58�;�^6�I�����,��11�b`9� sJ�K�d�8䬁(k��0)�?�	������$׶L����4��O��Z)K��n��s~bUIN#��.�<�UB:P���ʋ\F��n")��W����Jdb�e��Ϣ���C�֤��Pi����&�&�p\mX"*:����|�4���ߒ��]�6�i��h Wb2R��m#�"aiCL���T֯�"�#�ry8�?mH�1���c6���B�Xp1ޘT
c/���F�������q��L*:�H�=0�B���pn!c�8���.cC�:���q^<Lu�����h:���h1�d6�ԑ��~J����	�q�
��q1�&�?��;q�P�h�_ ��A�M�����JWkIɉ ������ܴ�D�_��rz�~�n���1��+�ԇ���x�)�TK���f��*2�jI���<BF����D��!>�m�{q6>��r��j����q�b�ɰr\�%d1�"5��q�N�)�&�������\b�[��V���P_��xY�LH:�+�%��3R�q�cjăk_���IR&և��=�>Y��΅�gC�ᵡ\wJ�5o��kBDĎ�mZ����_u5�c_W5�u6�
��*���tU��)RRZJ�)�^�m�H�4j|DB#k�������%6�fù��{H�+V4��&i ۷����F���LjTOm�KW[z�|,���A���vmU,�ֆ�Hy|"n���S[z0�חkMf�rS|5&�������^��6��w�MW��mj���6���mbA����H6�Q��֮5"H6�[i�cj���A�6�F�(����#�Djb��Q��;�F�(����#�Djb��Q��;�F�(����#�Djb��Q��;�F�(����#�Djb��Q��;�GtE���u�un�����wA�Y���:�7Q�Qf�;��,Յ�J���J���J���J���J���J���J���J�ƔƔƔƔcZ�kI��2�&SbL�ęY�YYYYY���� sK�,|Xic���YYYYYYYYYYYYYY	��K&�8M,p�X�4��ic��ę��1Re�$�T�e�3&YbL�^���xw�5�޼,ׇz��_��U|j��U�5Wƪ��_��U|j��U�5Wƪ��u��5�[H�X�)�S6�A���Bir�5H5�q��5"R����	�H����nf�{�|�֗���,K���WS^�"ު+Jɣ#��OTӚ���YR(N��%�뼡)ii-~�m�+�=�+,J/[Me�"I(;�DI��I��}$s"kʝ�'x؉���l�(�/�$�M��=~�1	�/��E�z���X�SIi�Č	6�Y=f�&���Mj{����p���`څޮ�t��h r�J�jĞ��98��&�\Ɏ�F"�j;�ڹ�,�4)4����Z\�ޞ)_�Edu1I��hP^F:�-�j
ƾ�6�f�f�-��wc��F��10҃�������K	D��5i�J4�3+Rk���`�'�[&���cz(��GUv.���lu9���TE�h�!D�*)�Gi���'+�sX��*g�-7�Ɯ��Oo��6�Wdt�Ƕ���S��N��z"t'vչR$M �"Ј�1ZM0;�Ӏ��D)uXNV�I@�;��
��]<c�4�����@|�7rvi��������ӭX�:��JW�ʿ_?δ��
�HR*�(4�R�i�O5���gZ� Cm֤��|L��F�	���S)A��u���mM&��M����i	�)��"z�jRo�6��MX��3n�q4��r��/�2��p��1��^)3���1�&�?��Ɛ��F�Z�cժ�t`����ޫ�b��OP&�^\�$"0i��MY;��Ҝ=bIt�C*�{.O&��u�hk$Z��$����c��A=�
KJ	>�FŴaY���0�����iN�+G&�(�V����{���p�SHY����ǁM*L�W��xw���f����^�x��j%�Z�@�Б6�,�օM�|MO6,�8� �sh��.�4�+(�����|i��Mv��ʑY]GJ��y�5Kvu�����e�5
&�%&���׀)��m��cd�F��B&�^��RU���r��V7Q��#�&ݾ<lo^ے�����;�&��H�W:ߒN�M�������#Z�S��)�+9�H/%�%"Ԁ��pN�my�cz�\tAj��sm�6�&ډ���H��F��5�����m�km#[iډ�A�km�_iډ�A�jD�6��k�#[Z�m#[Z�m#[Z�m#[Z�ik�֐6��mik�֐6��mik�֐6��mik�֐6��mik�֐6��mik�֐6��mj#SCSF�4��(�LiLQ����51�51DjcHjb��Ɛ����#SGtGtGtGtGtGtGtGtGtGtGtGtGtGtGtGt��J��&+LV�"�XV�
�aZ�4Ն*��_�2�'v8N���<H��O�e�/�,_X�,�|Yb����e����z��W��\w���qޮ;Ն���V6�V��Պ�UXڱXj���Skun���6�M��m���Q��6�Fۨ�un�m�m���[Q5�[Q5�[Q5�[i��㈬��;�-��of��
�K���eu7����Z������IX6��P#B��ڱDjM!),����*��r���;�&��"�'�Q���:)&%�`�N�RY6[Q���s��`MR�jvk[��.<
տ<��,_��%Pz��5�o&�m@��xCH��hg��������GW7Ɂ�bq ��Qڨ��e �E�#P�вR�JJ�YIL" )���N��eX�)��ti�`mo[�h�{uq�a��Șǜ��I���RkF,��V�����Y.Y�� �b$��9L׆nM/`���rמ5��VN+�UJ&��k�&��6��ڹ���T���;��Y��4a�����(斀��R���XVDW4�Ja��r�v�>V�^UP�8�^5mZ�A�4�22�¤���*cF�$+���h<����F����������ǝ�P}�Q��7!#R��5z���ƕ���v�
�^�&�
i�B4��l]zt�t$_� ���
GP�u�~	���M��D������V,����Č+��%u+�o.%a��p�j��x*'Y��Z�����yƄ`D\!���Z�4`pc���?������!U���s,ja�~f�?jN�~48��z8���;�����K�h8�'���!��M�7ɥ���8?�������u�w��&O17��|$Ly	�9���{�
�D�<fbl<DI��ڈĜ�&�
��b^�$\�ѱ�4m�� ~o���
l���ХF������LԹ�wD�'V���������y&5T�%�<F��f<5i��5^v$�,H�R���4�DjЦkkS�%�L�@��qޮ;�Ƥ����@���T���Z��ޮ;,�6�x�����2�4�ͨ�Z]jj�kF7-镙��&v(R�V�sH'jq�ޱj�V��j֮oS+V�a]N�Ok߉i��6���dxԤ�?�EU#uj�M+�M�ؠ��.+�+�Q�"��U��o�#Z�J֣�
͗Q�I�6/��'{��ѽ~,��M+=�b��.��+W^�D嶵ꨁN��u��Q�iк��yD�c�5q-�ҰoX�:V�Jկ�N���:\GK��q.#��t�Z�-{-{�j$��SHڮZ��,�E�c���Z�8��E�c���Z�8��խA"m�Z�&�խA"m�Z�&�խA"m�Z�&�խA"m�Z�&�խA"m�Z�&�խA"m�Z�&�խ�M��[H�kV��6֭m"m���-[V7��-[V7��-[V7��7��4��#j�Hڠ�6�4��#j�Hڠ�6�4��#j�Hڠ�6�4��#j�Hڠ�����������m!f�j"�DY���ޢ;Ն���_6�_6�_P_P_P_PV6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�V6�un�m�m���Q��6�Fۨ�Q5�[Q5�[Q5�[Q5�[Q5�[Q5�[Q5�[Q5�[H5�_H5�_H5�_H5�񯸚�$IW�ֆ��ś{n[��5!�*�SH��U�ʥ546�g���t#��xd���r�\VM46�v]�i*��.ۤ���a`b׍��hc�@ k����פ���k"72!7c kr��B���Y�SⰛ�ı[5'.$T�w���H��ީ!7��6/J����9'\��M��Cw�A�"�x�{�u�q˚yk����;�)�si)x5x� ԧ@�%�S^NwOF���Ɏ��Б�I�nޔ,DN��8�q<�H%�)HN�Rpe�Zy�o�+����d�&���sP�k|�jw.�5�M�BA�D�-!Ңkn�k�m��׍�x��-��j����f�,��L%6��%���jUq8�҉�54Vڤ�A����1�x�0�QS^�6��Ra�bRY/��
�Z"T�.�$-.�e��٦��&ZPnnnZD`H$�l�&-��Z���ҥ�F�x�O)��C��n1��K%�H�p�Nj&�mh 5;�%�O2P�[Y6t�Ͷ+�ܖY?vv-l6�7����xM�_�[��D�xg[i%<�?m-p�84�0p�(�8A�!S�_�ۀ�#V�Z��z-��yۈL��&8~!Q�p���BgP�!�@E��աq|��j�i��j�i�����j�:�	 *Ax����|�����|��ւ���.:���x�T�ǝf��Mk�i9�'��@+h������|"&�ڭ�76��4m@D"y%#�U&VO��V���@mF�D��x�usA�$1A����̓Z��j�4�;��������0�1�V8�ܝE���s�(��Y�W4�%I2iĘ�S������Zۭ���:�H�C��{R�L���f$�3R���ejmD�1.W�uX�:1�M1jޱjޱ�ޱ"עH�Z�i���b���.lo������9]�.ܷ�[��º��.�2l,�-BEJRcu�)�8���V�R�eR�-�}6&�8�Ϧ²q���p4���VG
�IA�Br�~R��Jm�6��K���SZeX�<�;�,��H��d#�4�$bLM:�Kf�8^(�ڜ67���o�
SQ�j�L��/�3�i��9�0�&֦��K�	�A5X&�T�+$I���`���`���`���`���`��GK��H��o���M#j��t���`t���Ұ:VJ��X+��ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ�ױ���Mm���Mm���Mm���&�D�H�im"m�M����6֭mj�֭mj�֭mj�֭mj�֭mj�֭mj�֭mj�֭mj���k���6���Ik�:��un�m�m��Z@�H���6����5\M����k�$�HX�6� mb@�ā��k�$�HX�6� mb@�ā���_o�x��ƾ�5�񯷍}�k��_o�x��ƾ�5�񯷍}�k��_o�x��ƾ�5�񯷍}�k�S�jt�N��ҵ:V�J��Z���j�+�ҭZ�ntb@�)�mE}q&ƾ�& i�Ed�e8���~i(�KI�@ҧ�ǭˡsx�~;)�&'0���NYp1,��E����ہ~�:'��mz�0IN~ZvY$
a���hU�շ��el��?:&'#�U��I����܉�����n��.��s5';�'��
?l���#Ze��t����Li�%�\��*�`oZ5�2�Hy�E���H��G��JV�NI6���0�"H8�M��Ԝ�koF?�i���5DB>4�WN��T�fbhX5�7��M#^�ս�[ډ����Q5���Wj�mx�׍�xj���Y��5]m�$�j��iA�M\�4��6��F�⑉���l�����5d`�-_��E"y�`�&#S�.�]Ty.��K�*G1���w�]���꟟�
M�2�'�7�&^C��Y�~�mD��#�St�����D�{!J	����74�u7�䢐�H�V{i����
f�jj�Y��{��e9��lQ�a�������|`DS%��
�)�J�o͡`�n�(.�x�uj�D��TJ9]J�H��B�D��W�2��8�#�E\�t�`�nu+�HI�0p����/��h���¹�8�բұ�?:�����8�#�A�u�#����j�i�|�ۀA||��P#�	O��|����))��z�<d��1�e�P�"x���4��h�n5#qK]aq�0I�z��N��"%ʎ �IU8�"J��$M[�3�Y��f��:
o��ú8�D��!m
S���*����nO����8R��]|S<�;�_i6��k��@ԩjS2KRT�R�ݺ�& 46��r�Ńj��mPi��{X,�&��7����Uqd�@ԕ Y2�mN)�G��D��!�z�Q=�Sz�o�,�QM�zd�8M
'�S����؄׆47��$JU�`��Z�mi�y�0������LNi�U���պZ�MI���۽Z�y��S,�7+&��|qL�\K �[PKR[eL5n��ճS��bn�����#c�ܻ�%J���j#����^Qᶂִ��N~�����}Z��U�ĤA�X�i�8��n���n�[v�۷�ݾ����o��}R��T�`ޱj֮iV��ک`ް֤�SU*j�MT���5R��T�J���,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�+{R��+{R��+{R��+{R��^�^�^�^�^�^�^�^ūZ�խAj֠�kPZ��-Z��jV��Z�խAj֠�kPZ��-Z��jV��kkV��kkV��k�$���rA�D�kQ$�HX�mi��6����5\M���f�)[V-[V7��$�Mᵉ�xmbA�D�X�5�-Z�Hנ�km#^�խ��z#^�xtcxtcxtcxtcxtcxtcxtcxtbս�[�ս�[�ս�[�ս���^�^������ă_H5�_H5��ҵ:V�J��q.#�`t���$ͦU�7��jx��LQ��U�k�b���q,�x�v?5��	�`�����:%H��A�Bo�B��X&�,ͮf$�ryY�mz�+$�7�QGGC�4��|ژ��V�����DFZ�!%�=�z�Э����#��[��r2���'�0-s0F�����h�ctzt�Q��y��d��h��@j� ���a�M��:��c���a@q5&�N�	�"�%�AО`�LT0��M� �۠�$�>
�{��O$q7����Dv6I�"��*�ތR�DF'6�蔜N M,�,O���r͵D�kX�oPH���z��Z��k�i��6�mm&�׍�ƪ�W��ʦ������)�V����Vʰ�DLp7[���b�(v0<jw�	��b�#l.]A3��r���-�9	/�Gf��ۑ��B	����F�Ɇ�21�ÎEҀ<�&~�VmPY:f�h�<Ԥ:5I����D�1�"��<�����ԇ��׵��c%��*l��(��S���f ���|��X��Z�������5h��Z���2�_���q����
���|�F����9�%@D`D\Q�p�q�����+@�HqQ�,�j�^��� �\k��q�Ƹ��/;q	���A(�������p��:��@��(��|�� �h8�ۚ�`Һ��ۺ�b&ݼQ:�+S;�Z)ƃ!��Cz�I����9	b�X��e!��:FnI�H�--�\��:S%�%b��r�û��ܷ�!Y1jt�M�Q�GF7�F:�O�$�DޞI�&�k�ѷ>V���d���c_u&�����r�ک�5G&�%r�wH&k'��MIHE�sA�ʕ�A"��ԕ2��R1`֜X��Bs��Ď�)�qQ͇C&��Q]b�X�4[�lD�GZ�V�h#�h H��N)�
�5K|�NR#�����e:%���T�����6�\���H�j�!�`��ڪ&�A�b�Ϗ���C^�w�JE��D��\S�S5��"�{z	�h���O͹��w�R��/���f�N$��2�Z�ܦ���7���|NPmS���+|��o��`���u:����۬��ʳY[��ܷ՚�۩+5��YT��L�V�V�SHڞH�Z��7+�4Śi�4���)SLR���M1J��SLR��T����5R��T�J���LY���M1`�1J�b�4Śi�4���)SLR��6��ok6��MT��J�ԭ�J�ԩ��5R��T�J����8��8��8��8��$Z�$Z�$Z�8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��$Z�&�D�H�i�	��������������k�&��kn&��kإkإkإkذ:VK��b��q7�X.&����ޱ`t���,�zŁ��oX�oX�MV	��5X&��`��U�j�MV	��5X&��`��U*i�c�
c�$�"i�&��MTM�D��}jt�SU*j۷՚i�c�
V�S������XmRy0�Ll�����R X����5|�Y�����ؓ��$�MS��kXo�$���Mm��{�p�~q"S045��"����j�_����A��-SQ�ܛ����7�`4�6�7[U��4�Fg/sw��_���̦��5;e=��%B�=�9ߥ�9 �U��5��*	Q���G7vT��A1��:{ۑ�z�5��)���Gra�L�~&�@��Y��@/�ңA>��9��7G�Ԇ""�Y��p6��j�R�&�oK-z��~(�"F��gĲY�ZYskM/b#�u�mϖ%�)H���'�����Ǔ�e����q\��)��4ěz�QыV��mkU�,�uZ�V����k����4�H@�d��ܴ� ���9�n�9��Ҍ<�uSB�\��(1q�GNPP~}젞�*j�#G^OV�kV��m�~�7Gf�8�-MRk#�ZT�Y��Ev��D�18J͇��$ޒ'-�J Q�2�ܲܓ��4���˛�pdr� N�3�x�U1Al��yLlV-��X�����r�`+S�Z�u��0�>f����aq�m������	�c�s,��f�?�η���-qhX8�p���N� 9n
2�
Ԃ��tW���(��&C���Gn!3Z/�(c�D�	�[�t�W���h�1��%<����W�d�0�RY���Ւh�K&��F��UT�e�C|,�.�sĖ�^�]Egz��ބ�q��i�A��Q����H� �<�O�I΀�e9�aX�ڕ�ڴJ���b���\j���G�f���o\F��ᵍ#^���AXtD�oP_7�_7�H&�#j�ݠ$[nR�3�ubmG;���
E�T�k�R���RrȺ�X�X,		i)=OnM r�z��nb(\�m[�Ѷ��ꔬ� �++���䩥�B���jS&�Tv��	LSlRG	�$�&��`�A�IMN�ɯ<DWj��q�9d�8�ج`�j? i>0+�6����<�@��oH$�:�Aem�Kj�M'��;�-�\D�Ok\��������bxؒ@쒷-�⺑ k��wCA��q,H�ɾsz���vbd�����n��Z�$[�,ӆ��"sz�_�MkC�cY�$������5*��X�б`�H��D�X�֧b�c;)*e�L������
f�Z�Z�Z��d�n�[u#u%�R1�RVk*�eY����lY0زcn�b�b��b�r�@زa�dŚ��5#��L���Saҥok�ۦ��}m��n�Mm���Mk$k$m�%+|�J�b��b��bE5H���J�����4ś{Y���ok4�m���Mi�����S[}5����kMVmkm|��ۓ�`t���Ұ:VJ��X+�`t���Ұ:VJ��X+�J��SU*j�MT���5R��T�J��SU*j�MT���5R��T�`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1`�1f�";&���V�E�bA��V�5H��ҥojT�J�T�)�d���\ko�+�v�и�޿,H&#Ku�WMM�b���iY6[���YS:*U#�^�[:7]���gCɨIe	)��Ԟ����cHV*V
o'�S���PS��)��E��SI�_((�Ӽ|�@Dd���$|��t4a�!�۵궁A�rя�Kh���O��`]�-�o��
U9���a$��b��˴Ě�
qև#+bj
M�"�"�D6�)�Z�j5�L"&�y9J6-T�-��5��a#B�LKn�T�I�k|��u�[ăjS!��F��h&7 mi5�$�T<���S��������ް��ho	�7m�)��(�V����U��s|�A�D�kؑmi�lSԩ��ԃ���sh5\�)?+��m�\��mO���4�6��!la�M6��%�Щ�
�Ar�c4.J\�t��=��si���-�5ZeRF��U�<1�G��4(-�	�@�av������ɫ'B���t[u�<EI$h$�&L�8e*rrsZ޵�3���Ltt���:D<`�w��M��S��ؑ�80 ,�Nz �0]|�e�i	�ͤ&�����t�@yӄ�Ȍ^��b��� �����T(ߠ�
�֤6��̣=��#,o��U�M�zC�~!1��a�-��n!��8�p����1��`�4���,����Q����B-M�:փ񈘥%�֫�sf�F5�b{�4S Y5�Zo�SSԜBS��d
��x�*)�() φ�N��AJnצ��Q=T1���	�`�aH�[5;��O��2L�x֪xߚBj9��Th5m��i2cL
k(X5��&�խA"ױ"tA ޠ�M1\��[T�&��'�5&6�&ܡNMO6�]�D��a�a]InZ��z���WY�O�u"�[|x�w O6�4���4a�ژbt?ېh�rן��V���H�~@"r&�D�����}'��)�y�ri�DNj��&���l6�w�&�ge�1�I��۔��E�j�H��V�Ԕ5)��F%J��W)�%gf��Gm��8�Կ~6���/�"�T�m[6�0��\I.��&<�$����I$p�.�oZm�e�M5����Nk߄JDB%����U3�htDMir�|��n^WƳX��(5eY���I0֧DOX�),W�+��tF�:#B��bòŇe�
�D
�D�D�D�"ʑ���5#jF,ԌY��R1f��++r��L+�6)m�(,(,�+���⺑��2ŋ5�ʑ�v�Wogf��MR)��eY��5��Y[�#�#�"�"��#Z�n�A�Y �YT�+���[��4��4��4��4��4��4��4��4�3}S7�3}S7�3}S7�3}S&���v:N����m�f��m�f��m�f��m�f��m�f��m�f��m�f��m�f�ԩ�)SLR���M1J�b�4�*i�T���)SLR���M1J�b�4�*i�T�v�۷�ݾ����o��}m��n�[v�۷�ݾ����o��}m��d��H��H��b�n�cn���V徕�SBjWo��}mԕ�ŋ�:��r@��iX�,�\�@�<��#��H�- ��	Asty�0H��%:�=Li"+�4:)�52�ܷ�����&	1L�WS�/�Ą�"yY��VI o@�5���i')Aw0�hɥOtH�.�X6�<ho��M��׷�%��$�ͨ�Nݟ%{��_G�PF��� Ҧ#�[
�I�:��L8�/=�\�`䎘��6�D׉�7ɅF��3i���Ű7��i�H�~f�\`t()�GB�h��1���k: Z����rkz��&��$�'�IP�ݽ)-���+z�<iR&��Gp�V��i%,��#r�\�O0%��M'DJͽ�[�-SH8�H-[ڱ���x�TGDK�jk&����xiGH�Vےx롽L*Y�E��V�ta�v��%\q*�ǐ\��X�"T��`��9=�[{��A�+�i�#wf9>����#[jB�9[)S����"�D��_��b"�9�i���p%�L�r��zޅ���v�tt��~�"p����ܗ�n�RѴ��x������n!��c�è�F8A��!SZ�а�za��Z�u��6�u���>q�r�`+S�!���8���Хiw�GW?��hD\�0�M�#�b���Q(�"��V:�us�Z����GH� �6�ܤ_
T��^7��
kZ�	��d�ۅەa]`�6�J�U!��yd ����y$��GA�u�o��E'�]�*pw�7A5V�K2���A��41���P�� 	��;����jtK��*��Ь54�IIq_����aY�Xi�k�R��R��)Z�m��z��4�E5V5�5�ҿ���Гt��$%��ӱ�u&LQ6�N�*ͽ�SFR'w"y5�� �VFZF�ɱ4�Y^�[��L�֧�����AsIX��4�N��$vԲ�X�Hͪ!䓁��ނ&��&��<�&�'5I�V��'	�JDr�0���kG[u#�0�����ײ�`�&�tvl�����Hj�S�\+"�;j�6J�Ƒ�Q��	H:�� <VX��Z�%�R�z\�ޗ&$�\���k|�y#�H� ��/�?�0hS��
Ά�V�%Z��P:��q5�M��N�����)�O!)!u��IR.�n�Ew ��]N���DlI S�BX�S�S�S�S�OS�OS�WS��y�O6)�e��)�52ƦX��I�I4)&���,��Y�ئS�;)��(��Ge������Wo��}Z��U��Y[���R0زa�d�bɆ�"u"�"�"œ�#k*�em�U��ko�f��o�f��o�f��o�f�lYM�)�e6,�Ŕز�Sc}nN�1�v:N�|֚��SZjkMMi��55����֚��SZjkMMi��55����f���U�ʳYVk*�eY��5�f���U�ʳYVk*�eY��5�f���U���5�f�b�eY��YVjF,�U���5�f�b�eY�ܩvX�L�DkS�f�b�c5�&�����Ԑ���X�k�N�*I�Ј��Dܝ�7�v��gG3�ؑ�uHֻ�;%l��/ϓ�4ϑ7��B%��\Ha]ꕹy4)���$M�jd�m5z�#ȍ�j{Z&���'�F�6��Ee����hm(��9���T��ֻ��-Q��R�$���y�|�}v �l'@���M*9���(�d�d��Y^�z��&�4���1�U���ų(=��F f�3�zb�mm>s$��˓���rh�R�[��PH�17H�O%Au����В~_���%w bB�ja!L�j�R)�i"i��mtk^G���p�@DLP�� ҹȲ�|�T�&�
� �\D�RoPS7�6�$�$��$�j�M\)���e�ڜu&��)+������.k+6��qS�:��x��TY:"j�h�A���Td�ǐ\��1��AR'�� Knkm���jc�u8R{�qQ���H�Ғn���kHܐZ�i����	���A�ۀ��oGF�''�\��Bi�
MW� �%��p�Odh�i0�L-7j�Ϛi�A�݅{G���޷��� �5��@�۫BJg�Г&���c���;6�Һ��۫RƦ�x��w��u��V��S,����ĢQ�ͺ��kF��±1�4��=xlR�v�"�Z���gXIL�S,����j�:�N�j�:�N��"���O:� CZ����q^#uc����gR�
�#�=�^HK2{n�6�J�S�ȏ�B#���$�Y7M�'�\�$ڷš#A�m�z�
CU�2�T�OB�"\����1��2�w��T�fѹ,J�,����J#Q��WI[��ʸ��mE-M�[s�s����7)����m��IV	�ƃ�AM�<֚��R�L�O-	���Z�ܩ+�J�a�NpD޽�]�
W���=b�LX��
Cn�b4���y%6�ϖ-�a��$���� I��ޤ^�����L-Y=F���E�;H*px�L�_[+���b��S��A�W6���p�V#�r�m��6�h�s�հ���޹)ɡ՛�x��#)���=H�׫�5���.iz�Kw�I.!,R���!8�l����}����O}R9���㺐�1��Z�Sx�%Z�$W�
ƽ�&5l,�d%���a�%',b$�n�$^LY��;:�$�4:4:$�NS���aIN��pA�5�'�$�����b�WS��y=c'�d������2z�WS�i)�%+��	)�!,P��	$�u<����3��kRV�{x��ԓ��vRN�I�I4)&��,4,XhRN�I�I;)*e�L��Sb�lY0ز�L6,�œ�)�d�b�lY0ز�L6,�œ�)�5Y��彛ٱe6,�Ŕز�Sb�lYM�)�e6,�Ŕز�Sb�lYM�*�cS,je�L���52ƦX���cS,je�L���52ƦX���cS,je���b�2ƦX�L���,S,je���b�2ƦX�L�a���C��g�pVnr���SB�pI�	���bI��IЈ��@��`��J���MU�L�ɻ#vp5]��i�bM6��TiR��l$�~4�a'@��]�	$�$׌)�C�"5sz�ځ����G���j�ց�5/ߚ�;L��n^����btQ��Ev��c,؍\x�|� ����	��/ٜ��j�iF<���ir��$�h<V*J֘[)g&T9�9''�,JRs��Bz�5�k|�����MV�����[�g��Ϛ���:N6���� ��4��t%�45���dS/ϒM��hӹQ�XV_/���h�RDH,�-�2��4���� ]��w�O�J��%��.�'��)RH�
uͺ��d��eH,����S�E"	�R]e�Ij9��{6�F�2Н�-��ƫN]-��auFN"T���Q1��b����1�QQP��~�&�;������`��JъE;U�t4�ɢ����RR��Nα�Ԛ�h+6
�L��mR����U�Q(�I�M���PrF�&4ӈ�L���R�0���F��x?m-(�k�q�1ša���Ë�
�����?���0�p:ޅ���J;i��M<V����qhX�Ƈ�m)��>���Z���Sa�Rw[��JQ�H��@�L:��&�u�и�+����ܯړJ8����p��W�H|?>p�m!F�-@p�a��u��Cp�e�
V4�'�&�v�$���f��iѯj��S�E�yI`O,��֚%J���*�͡T���M���X�7�o�A$B$��c^xв�
��1��J�6�Z��%��*�4łj�7�Z�5��+��hY WY0��[�����%M,O,�����3�~���+}X&�����\RS��[�a!��9=�n��NcU:y��`tw�oN��⑹Mf�;��V�N�)��Z���F8A��xBP�I��_�'D�8ꢛ��5��4�&��n�6yl�~$�$����?m�ƲF���nW�d�6�Il��H<lp[�	��`0	�e�`
oW��]�p��2z�	8��j����
��K�0A��%J6���r"+��""ɩ��=��!:��ޭ
g;nֻSO�"��	<����.���n]�B�Ry0��`I	/�'D�蓝��"yDO(]��!wD.脞P��hp0$���Pj�S�Jx�O)�$��)�S8I0D�a9N��w��4$�$�ا�U�JlS��y=O'���<$���0��X�KIc'�d�$���Ԓz�hRM
I�b�B�hX�Ф�,4)&��
I�b�B�hX�Ф�,;,Xܤ�5���-ʐ��I;)'e$줝����vRN�I�I;)'e$줝����vRN�I�O6)��<ا��b�lS͊y�O6)��<ا��b�lS͊y�%;$�d�쒝�S�JvIN�)�%;$�d�쒝�S�JvIM	(I$��I�d��p[��pT�	�%;�w|п��N�E%�#K������D�����i�1$�sM;����"�d�k�CK[�l�0�P�ꈄ�JSt0�74�N��)#���b���N�⑩�BkS��9��>��A�ɦ�4���˽������dH�D�:(���j�;v6� �n��ȉ�1��;�v�K�_9��o�RO�e$�K"hG)�*R&4�{*[n�5A�9��;���i9N֒ޮB4��y���EG�S�T X��@ȍ%�ri�dD~5!7HE$�|��'4���|�58�����y1q���m��D��^ږ��V��D<wH�	j潯!	�7���U�L#l�����ٯp'�6�%�W�I�b�bʰY[�%�_�E�%�����Li+d�@bk^~�H��Ԅj��o�c��H��Mڭ �D��"�� ��r
�1rnN��eM��d����li����N56��RLl�"r.e�+e�p�ב�%a�I0�D�?S$�\$櫈��v+�J���Ǉ��h;�hi+����O!&�b��i�{�p��i���J��@��y��pBd6�+�� �jj�Y��|+�Z�ZQ$ۋ��u�V���&�RƦ�+�C�D��ZG�`����ТI�i���Q(�����I��|c+f:��c����B4$�Jg�r�%h�h��;:�J%"�n���7����VR*�*A&��� �:�v��vX<T�cx���#��"8�W�2hIĤ;����!#�ޏ)�i&�1ޱPN72���bo��"sdݫ˪hhbCCU-0rw���M�+7�� ih�H���A|Rs!�/s��Ԏ۬P+�&�ҥ3}m��x�cx�Af�@бD"R")����dx��h)���D�ִ���[��}f�cr���ԅ�K����iG1	>�	��kzn&~���l�W�Ƥ��k��׃GG��ț�8�#�^�o�BD��X�Y#t#^��Պ���/ѣ@h�v�8��?��()�,���D�q7����u�R�1"$��<��Q�a!�|M,��@��{�t�lSaN�p5����H&�V.�16IoUF'�ᩩ��Nn�N���a6���t9�4Gȋ� :]���Z�}t$�7��mD�,��1$��\�!�'�s�H��JKw�Bw��(�;=f�����]�Z�5_�K��&<������B_�K��/�'��W�tDN���):$�������yN�)��:$����\�tA�]�!8 ԓ��	$�I0$�`5O���<��T�j�S��x5O�`Ռ��T�j�IBI(I%	$�$�$���Rz�OS��y=O'���<����H�n����j�Q-4 ����2z�OX��y=c'��������2z�OX��y=c'���<В�SC������a�%48hIMSC������a�%48hp0���{�OtI�=�'�$�D���{�OtI�=�'�$�D��T�BJvIN��48I0�%!	I�Y=~��TLz�,�N�Ӹ��R�k[�yL�$ڟ����F��Cz@���.lS�����ꉊs����6ڻ�7���E����S��0lu��Hp��",����$��V �b� o�cn@� �ܔ�e��T�<��RSy�Q5�4�v n�(PT�?=��OL7l�{KK��o����i�w"<�GZځ�֤�����rT�P��?-R���{uA���X�;��7[ :|&Yt;���4��mNy:<�8���'`�B�f�oC��L��>_��thٴM��D�x��4Oy5�#�h�l2�٦�M��~��%�:	�c�����b���8v_�7.���"z��Ք줚�4��r��]`�J�,��
�KR�a5N�B,�7&���đrp"B*9���O���Z�cB�"T��q�H� ��a�ɲ��-Lkƭ�� ۘ���5���L6�Imz4ڧ7w�	��MD�!]dމ����MiB�4��&�R��@jFމ����͆�)8�LPOsn�ݍϓ�#�rv}{ ��P05���``���n��n�)�к@�"uM��ZDrvmդ���l��J:��y�iʙ`�n\D��Ԇ۷���J;6�ӳn�Q$ۊM4��`����D�n)Spp��4`�>!�@EhD\_<G���_� �I�րV���%��[C��^�0q��0��> ���?��*����?�@S�7�Fi/9ܚ~ ~�#M,�RJs�Qd��1��m2�"�d��7j���2��P�.�e�~��i�#j��MU��x�VrnIͅ�٪�!4�F���2kR*��M.��+���X��p"Y��H��%ĵ:�s�Lt Np",�N��e�Ԙ�t,��M� h���Dw�N�F������N &��i'z`5LY+�EH�Б�d֛Ze����\tS�\�Gt�:<��J4m��16����A���%���@7cJi<�tr57����\�`�)�Vm��T�nZԚC�� ��V��OLn]��ے/��2���2�j[X�-�ѫ&�d׈�
G7x�Wx���ȞD�4�ߛ�e���S���?*JFD(��aj��F���� 5F����^�M6��D�
�J�OQ��a�긚�a�~��� 6�� 6���b_�OY	�)=e'�$����"w���5����|.��Q�"tJN�9�'8$�D��SB�h_�O)9�&�$�D�����My0��a�$��и��@D�D"I p I0�`5$�j�S��(]%!)�%<������BS��(]��!w.�����pA�&RL��I0�`5$�jI�e:%�z��6�;�*�Z`I$��JI0$���L	$�$�I(I$��JI0$���L	$�$�I&�L	$�hp0$�a����I��I&	$�hp0$�a����I���{�Oy0���L'�$��	�=��{�Oy0���L'�$���5O��$�$��RL$�NI NI b �D�'�"{�P5�x��S DbF���Id�z�:;�	�R����z�S�D��^�t;����'��"6jR
X�[T���$qN�<�)T�Ge��g�4a�t�ިV �H�Ky��9�P	d&1�~	~�{#~OGl.F�y	�->}������H���7����C|D@�KR�(�t�c��2�Sց�YRQ�ˉ��\����^�)5I�e�����sL}~?}i���DbD҇Aݺ$\m���B��Bid)��TiS�-DN��4s��)��G�#�|�6,�gC�u����瓴H1��u���zn�&�Js��Hj	���{�j�8Rt4�K�K��b�2ŉ�*E4dH��ixRF��d	�Mf�7)Y�ԀkV��� �KT�͔M�h8yq�A��{G<(���a��<����ש�Ph�1Ce�x���IS��bفsI�ށ��@��F$jE4�Vϛt�a"w#Y�j�Gk\��֭6��ƚq��{T���@F6FDZ�%���0����p��0�D�1�$��~|�����z�=�p�gPGn!0��;�!`ԃ�q�m��t@7������6�y����
��>Q�������8���;���ҫ��4���F^����ڿ`V�ZZ�9px��r��0"�u���@�J�����:������/��,�L��n�Cbg��L�މ��Dk�T�A@�A��>S�M��.Щwf�v��on@�6O�����!5J�w��Ju�́fھ��wz#B�)	4p�ڌ17�[��(��%�wແ���<bI*1:V'�jD����QH��+�=T���V�q$�T5�Ĥ��9M4��5��s���*%��Au�$St+[���" X�����{j�HF�Ĥi���e4``&�,��I�i9HS&�ִ��SF����5M���ޣ����Lly6��Ӻ@��Z�8\a(��u��#s���Xj(x����U���ս jK��BZ;xޖ��+��d��HP�r_�k�V���NhF��rE���N"%�����F"����6����X�9�"7�۳hڥ ��j�kK'ͩAu�u�Dq4� ׽Z�z�;�sz�@��\�'�	�V��;���|�Յ'�BH�w���w���w�	/�_�$�`��/�%����R[�KyIo)1�!/��|�[�5yIo)	!;�U���D޸)�I#�k�P�䨘�\Lt Bp0��`]��!t�D����RIJI)I�'8%'�������w.�`]��pA��&\RL���p VS�6������.Z�6��Q�"yDN���:"'�D舞Q�"yDN���:"'�D�Q�yDO(]�<�w�D��Q�yDO(]�<�w�.��P��_�.�����u��(]~���_�.�����u��)	';�09�b_�*vSG�m�v�ރ��WR
).+MS#R���1�j�ɧ#h���h��_$��CU�IM7�$����NQy.#J�N��qAq�u$�T�z�4��ֵd�� {j�G�Z�V�`h�)'����ۚ*=�>Z��iz��YA܁��1٪\����1�Z��v-{}O<y�r�K�kd��i"*rS�ܑ L�Ӕ
��I舃#�(\D"3RI��"m]�^�;�ӗ��R�N��Mf�6�����)���.~0{1+�guq�9~�א��ƭiieH	�GRo��ԂO� 5�'{a��F�SI	�&�	�{Ĥ�^F�m�d�@�i#&/�&â���*I�� D0��ڸ�D��4DZv)���W}J֣�Z�rx�X��G
�"�בŨ�uLL 1�v�
V���;j�p��t��N�h26:P�R�P�����%D�����1�|�_��Om7dB��!%�L��;�čz��x�m�@]|�6^�%9�I�D@ �t-R8�&�rj),KJ�́�#O��$ܷV�n`�ϓ������S�۪��0ZW8G�A�)R7Z�~V<Le��GV:�w;�I��S��Z�����i�20rF8A�oBM7����p�i�S5�G*$�qR��:� H����jCm���� ;6��ݼ��#��Ԇ�H[v�"�X-iˉD���η�GZ��ݼ� �����W_(�-��H�Vm���x��G�A�S-^"%3��Q<SFӸ�"�J_�n�Ad�j�$����#��MziA��C2Ш��2�h�s �R� ��|`�qJgzɾvk� �G��@%����q9�{1AM���m�t[R54(�<�2��� �w�&����!��^���T�C�-���y��XzYz��A�ש��^�6?�D��xiZ���SH�^~ړĔ�r�y�C^����5)����o��'���ې�	�u��
Б�r"Y6�WAء4>!�ͪq�#z�x��H~MOz�+�V���+�6�+z�p�H�y��N�sJh ���)��=r��b�MA�w���;,��<�HӢ��~"F���"��`:�vt6��5;����w�]���U�z�oG��47�g�|?T@� 0<�_���"_���U0���К�%��؉Hq�����jI+I�TOV��ɠ��8JL�W��#-���Iވ�I)	J@r`�%�cW�j��^���Mw�OX]�)=d�|���S���9ŋz(������bp��8jF�oT�t��|���RL&���8"'������RtI��9&/�ǔ��aI�)<�RtJO&�!:$�!:):$�|����E�)����cZtBw�K�	�!/�'|������Bw�K�	�!/�'|������"_�D��<�%�O(�~��Bw�K�	�!/�'|������"w�N���;�'|D��"w�N���;�'|D��Nw��y�4�.�h)��׽k*�J֯����f�Ȥ�Y#@��G,�%X�1~oI�T�f��c������mѢd���<³|�ֶRN"07҇z��9�;�MM�z4v�y#��Ҧ�v��n~�?\HF0LL�L��a�(L5���m���а)��M���M�9*8(6 r}�R�tw"�t.ieNQ���L�6�%�_\���%����r\��(�#�7rz���ɢ2ҲI�L;�J�zI L')ڦ'�H��NP~~G@L�A~|�k[�at��'?ɊBsԲiF��6��$m��j��g��ܶ�u���M5�DI2��Lt-[P7���m*Aޜ�mL4��
�I�ˣ��l�L�V��R"y��I#�u�	oX��O���X7���%Ɨ��k��\�Z�I4��v��l�B�ci8Ҡ:QE�<)��9���R8K\��"Tqr䨐hb ���Z~ZHT옶`@P�:$��DF���j�$�t;݀�.��&��uZ�ĦoZ�h���m�`a#i�HZ$P��}�z��M��yО��9ͪ���N{"?l��ީ&�z�.I��d�H�i˩�c/����� �M|��Ʀ�Q(�5�f�!���E"�n	�SQ$ۋ�D��."Q�J�n\D��Ԇ6?�Ewr�%-U�S�D���J:��y�Jg��"9Y�Hk�"�n�x;6��2�h�iu�@
�zoS�x�;�
88U��H�:��­��8���N���V�5��hvq:ԫ塭&�#p;ۃhV���K$���I<�5S��'&'5��jce����.A�&B�cA曰�v�!����Db';�Ʀ�0�ި�֙�jn�X:E�ȁЈ��5�^A"y�Z�T5M���hI~�jM?�m��j�wkA8�M�ٴ�|�I6�D@j�����Tbp%mG���nD"y�4N;���eN�19:m���jkX���ez���H�o[+�`��9bm X����ĄŉSZD�Y4���7����X���Jw�����ڧi�����t�Xt1]ލ^K����Hڝ����Wz��Gʋ)�&[�b��L��!$�ב�D�(r �\�NR8LE��vR8LN��x�n�<���Po�(��#r�m�y#��'ᴓؑ�~:"$ <Z\��bڟ��"�{�Կ+-��͍��=H(��h;\�pFà`����Д��\j ��������_�%�J�r�D�DlX�)	JBR`�%��oY,5�]�)��Rz������s�Mw���HJhX�m�ɀ���r?���jH$T�%��
�d��-�\��JVz�`r��%�D���"tJN�I�):%'�	��5�';������L)<�Ny0����Ʉ�
O&�L&/��|.�@.�a-���I��	��9��s�Nz���';��	��9��s�Nz���';��z����@�����c�b�Nz���';��	��9��sՅ'�
OV��)=XRz���aI�Յ'�
OV��)=XRz���aI��BpJN	9%��P9��'��CzF�ZH�N&�o2�oS��&C
���:
�k���,��
��x�n�kڮ�Q "����S�d�D�&������	
̹'�ݮNt�ĥDA����|`�F��-��EU:�rw�I(,J�W�	헵C(�fg��E'��G�eHEg2�"D�H��R��*b[��Mt&=O����A�A6��jڢ'3u8��e�wt9��ʛW���tOi���
rlK@H��Oa'�Hmm�N�a!��޹���%������LZ�J��k�A�1$�bFiSt�:��;I�#��d	[�s�����|�n1̴Rb����nim�+#�L�h&$��"U2�����Y?/
͂z�Q5��Kk�d��d�I��0�vie6�$��1��"��(d��9�IT��W%D��41����	�<&˘�~D�A���U@�п#p:bDB�	ŗ�D�;6��a��V��F�
Ԥ"&5��ʆ� �Y���vl6+�"��������曛L�KnZD�E�u6����֪;r��IB�q�ik��q�_8Pq|�@�>��~�&8�,W�C�8���hq� F��������áWL���y���<ҋq���Ǥ7�h\k��zc�J��Jm_�3~>q�9�J;ip��ʎ��uqhX8�p���OʿV?ڛ���e�<oMX�1�*����V�H�Bp�=N�"S�#@ϗ�&�Qh�4� �ҁ�d�~�l��D�.A��Ar�L<�sE��dE����2E����)��a�,j:ܕ�!�PԬ�'���Mx�И_�D����\�ڧΎOTj�:�m���F��ē��|��$@ԍ��Y$�F䵊��ȹ8y+^&\�SS�)X���h��	Z���	�wZT�l�F��Gr������ �r�u�`�~L"O*?P*2�r��F&�H�ց�ׁ�-�&_D���DI�� �Hھ��Һ@)��I�T��<�]��cV�!��5TI��vO1�VN�A�m��6,�%wy�����KC���l�~~7}6�D7s;��$�E�#DK�F����mi�)������a�0��LX�ě���m �&51H�FTU4����򉱵};�T�k���KM mV#�BV�ꩽ��L_�&/�HV#��d�	0I��&�L��K�Ę5a��'��&�oY-�%�d���=:@�*D��f<bW7Ɣa��c�k7�-4�֏4^IF������c�I�ByHK�	&<�������@�7{	�V��%����%�������X�Sw���@j�@��@�������w�K�,I��9,I��9,I��9,I��9,I��9,I��9,I��9,I��99��sՄ�	�V��'=XNz���a,K���9,K���90L��L��L��L��L��L��L��K��HD��9Y);�O#%1�A6$����Dm���r�m�u�^�J�Ti=�o�4k�`my:�G�V�d�d�'�[rɈސ)ʓ��̍�er��9�i���M�L�����J�F�(w�<���g�� 6@���zhmA�h�5T9�OLG#[��vTdΊx3E��m��`�T)�`)�<���"��S��֩	�6��t�,��=���F�Z	��A 2sZ�$��l�?2�~��~niX���FO=�N"i�N�`��
����6��J	��2Bp�h���1 �œz~ם��I$ŒH���y�z�K-x�zm"S�'�/���t��u�ӍiB��0���Nn�sl�r*~hr���;�Z6��	M�TF�6�x�Cr� 5w�5/ߊ�y�0��mM+����RSF�i,��oE"Y��?_�̞�<��LbUVhh�41�*8�ȣ��	�T�`@P�o\k�G����yNY;��G���m3�S^e�E7}n�ʎ���|�05)��)�L�׹6T	ge3p�x���rב!�dx���9��F��E%+�?> ����u�MkD���%(��j`@r����Ј�C:����z���[�����w��zn�h��zkǀ�x/S�����1���1��8��;�p��7Z�ZQ$ۊ�Xu:�'[��բ�H�1��W�]fkH�ZEsSW:�媰�+��ۗ)"�ne*0�Nq6�3Z���$�s[x�S$Q��Ahhm�mx]J|V'<�7�kU�%;zH�kG��E��1��Zڴ�ӗX�r�&W!T�D�CPr{0Lr �Bn�#�.cζ�`Y)���#BI4֟��Iƃ[Ȧ"$Y%_�FJI��a�$(��R��]H�Yp?6����F��
���^�&$���׫$iұ\NX�)*;��M,D�)5�d�M�KmM/1�ryдx�Y6�iCZZRm��I�S+JC����٨�֘��i�����Mi!v�����P��hM* 8<�n�Ƴj��K*R����b��w?}k�g�$j�0�+j�l)����<�H(��׶"A���d�{��&�T�����܇
�k��&�kϒ	���D:(��X�Ώ$����`T(z��A���W��'�؀�n�hJi-l�LQ15�d���X:����e��A�I�l�H����dIJ�1�p��bY
kԂ��8ƽ�e�\m$�Q�Ȓ���s���I6�I��G���4zN�G���LJw�D�1)4JM���094JvX�)8���#D�5VOf���i��֤F�iR��1��DSR=��W"b�QM䈚�r�N_���9�'=XN@��@�³�VaY�)�P)��5w���4�M sH��+���`�ވ��@����z�_�c�ĥ1�
bR��1)Ly���<�LJS@�%)� S�ǐ)�F�l��j���l��j��
bR���%)�JbR���%)�I��h��<�4zM@�=&� M�G�&�I��G���	��h��餂S���K�'x!���w�-�:���_���H�[���8H���1�r4��Nj���:��S�bb@�w�\�΀Ƀ�� �z�#k�EF$����H��YS^�dґ�M	�Ԋ�E�mV����$1���>YɭՐ��a���l1�����`  Tx�=��Aȩ�<��$}##�l�^x����`ғ^�ڼ��8�������4ú���z��AP7���4��_�D������h���Mؠ�ו,�"�����ز$�@C�p5���Hb7>(TP6(L��$�S�
�� m^F�G���m@lI�n�n�<�-�H��\Lz�J漣v���t(  [I<���7A4��*.ޔ4�������!$�M'x�h�q����l�R��5�5�M �JȬږ�ǔ��Sx�V�&���!�{Ո��Z��CCEb�Q� ����<(�L��~:n�"Lj��)���LHS+5�j#���'|�>�	��R��&�H�޽Im���m�~�u�խ��Ԝ��\1t��98��m1���c�X�RX-^'SΦi����RS>G��_<���y�v�"ܸ�Gf�ZlR��)L�Z���=xN���`4��,�R-i�fS)$F��0$�	)�$�j��O^�β�=x;:�����_5�%����M���Ԇ�Z����n�RƦhnA�"��QM��rkH�TI6��/��n���j'h|C��>yۋi�8T"�ڑ�X�!�AMZ�mSO��f\�6H�χ������:i�3��=\���H2�$!�<�i�[r8&T�����nR'��ӛ$Cޠ�F����m_�<�뇉&��<�Fj�F�B��B��G2c|�Bp>����{�25t?���]$ �G)�P;�W5���z�Q�%��L_��4��bp�Z�l�����8ԍٯt"s��Q�uaL����%'ShQ,��y1�'�VF֐�M	)@om�ٖ��񨑠�ר��)
�#J���Q���j�R�ӂ�W�h����ۼ�����6��dֿLn$h�ۨ:��%c�M�a�w*}R�
�
���N|�'e "Du8]ާ;$����I�H�TM0I���"Ւ�z�R',Q����{^�tѦ�y�����n���Q'����ؚ[Y �̿8����MiT$�.֣fѹ�y�Sz�ht	"y ����R�^�א"X�[≨m�W�A-~��6�X��b�5 aX��b�Y@�%)�I�SH�4��bV��V\ּ����*:9/�o%"�Աq7��e��~p	17�`�`j�~kG�ѹY��cW�j��j���"��#H��)dI@h�@l4�W^���D�q�ǧq�D����[�]ވ$�`]ވD�DV aX��b�V aX��b�V aX��b�V aX��b�V aXzV���a�XzV���a�XzV���a�XzV���RH5 `ԁ�RH5 `ԁ�RH5 `ԁ�RH5 `ԁ��l��TR_�1*R5o&�� jX�,]�i&�TcU~�l���Œ7ҺIQ8zHה?���qJ�j������jDh���HK6�,�葥� F��VM!9���M�vY	�
E ����s�j�4
tߡ����%�0I��q����uR`i�@j{`3��c����'�n�%?l��"Zn02=)������T�L*Ol9#Zc ���w�*i�lA=*b���lL��DF�nYo�ͫ)�L�vN;,V���"r��KY�[V�hMNhp	H�KV���	$֖�8+�L�Vt�:7�й-HV6�,�MU;���R�4����VEF�u��9����h۲�eQ�T�jג6�ּ��m(8"8�;��[Wbp��@��׶	n�й�ܜi$1ޭiM�ܺ��R�H�R&�DB!�fm������Z6��%G.���*�hh��� ����-��Tu��m0F�EG�EIĆ
r�\L�bz�����Ju;�|�L4�����.mt)�����ԉ��1�M5��� rs�x�@AB�M�|Z��"�Hc�+�Y��sZ���F0I"���M�"�1�o���C���1���[��m���Bm����0p5�@yӾB2���!P+S�1��&�Z��t��ɶ�]00B�Bo��|�e�R���BC:��V�1š`��6ϐ��Ѐ�94��|�V�;i;J8(Ͱ|�/@����L\
(�[�� �_��i];��,QQ�-�!�#`�|L&��/�Wy-JL"k���B��0J��ED�
憊YTy�6��kUب�4Mɵ5�EM�0FU�3��Z5"4�H�ѫ�+�h�&���wPmHDJBihz��w�lZ҅F�ҁ1�� <KX�4�YN䓸�����hi��zͨ�-H��M/�Mh,�\x����bk�Ȳ� wy#A�q�Ĥy�m�9<���z��ב�N�z�ēK��9�w07Aok^�]���� �9 �9��^F&Sw�6�@�DoJs��vW)�/#t����b}u5���Wל��`�@jn�~���1�����4`�R#MG�{l��6��)=A#��M��j�Z*E�˽�c[s��f	^D��A��$TkIkO�:��n&���q���L2׹��	%+/�5�v��ޣgBI�m�����$��:��`O&��M��✎���&����Yadni�F摹�nY�ǘwaXzV�Ħ�)�Jw��(�בĒ5����P�<y�X�M�$�H����̦��OUJBI�Jw���!)�zV a���"�ǘwa�y��$"H������^G���E�$DQ�<�"��h��%&�JbR��#l,���6���#l,���6���#l,���6���#l,���7+0�@±
�+0�@±
�4��#sH��74��#sH��7)��cr�ܦ7)��cr�ܦ7)��cr�ܦ7)��cr�ܚI%�XK$DYF�X�� (DH$��kL���N|�&��&��~)+U���-~���58�ڂ9Б�h:JD��p&RM��iR��4@�!7JM�[���y��.����>*+	&7�ɋ#�r7����� 4�΃׽@���U�6|�P�`�$}7����n�L#Pl	�.v<�mS��:r���*8|���{A�v�\`�n�>(i�K}PTH�vv8)�p�v~�rG� 	��`�j�$~$�\���P�w�9$�^�H���d�Q��vkV��6�ipRN[��H��!	#N��CH�ɽ#X����yC���w*I8"My��֐��"14M5�S����S�e��D�5�JsQ��@�?mM��i�d����8Nt45�V�NKw�;��N�$Ƶ�k��`k"BZ���,���i4"���䛁bމ��.a�ց�E.hha�%D���*Р�8�y��8 �q�a~޼��sj׺ �����vz���[�b�4�����iY��F�"cz(�3�c�zb������SRJnm֪a�U$�_����	����Dc�2z�q[JѸ�WhI�DjEwSS6(��n�n/��u��Z��_�7��Sa�&٩D``�/����Ƹ~�!��]0�^���t@(���t���tp5�и��а�u �L:9n
1�6��F?��x����8�,����Q��;in#�xZmLq
���&JnB��u����h��'P�1�I(�@��j2Ex�Q�'�py,T��o�y	��rBs^�6��sP�4p`�(1��1rPХ.���Ss�D�F1���wt6���bhj�o��&��N�Bk[�ѵ�w����Gy�1�Tl�PPר;΍�#�3zHp�ڦ,ƥ
b�nh,��r��&�JV)�����ԓ@4�Nt�BF��<�|KkTMjpI�O&�KT�#�֭Y���t+��$�ŋ|Kk�R���L�V8LwQѵj���c�zH�qBU"p�=в_�OA���K}4;��d�����6��z�$�'|�w�!	^__�
$�T�N~�*'x"�aݺ�&�IeǑ�M�Q��p(>����ѫf�6�^�v[}�( ZD �I��|DK[''����;��bw�����:�oTf&�a�i�;���U�B�Jw�X�km����^Hƴ�qduQܑ��_�kԂ�-���d�tw�Y�4���mF�ja�m���F�YadnY�F呹��i ���h������m$Y4[V�ОtZ����rɰ�`�����p;�$T�$c�m]���q)�zw��w @�6��@���wa�y�q�D�,� Y@����.Mt%4�Wǘڍ�DȒ 4Ea�Xzb�����mF�5��H�����FF�Yadm�����jcj6ƴ����#sH��74��#r�ܲ7,��#sH��74��#r�ܲ7,��#sHܦH�HܦH�HܦH�HܦH�HܦH�HܦH�HܦH�i#	ò��H�iS��M%M�Xt�d~�@昒j�*�l�[<q�1ډ;=[� (#[	������0�ږ�K(�h�Bi�S��GS��"��6�p����״�I�#�����ֻ���E')��0�`�$��TD׿)ȭ���ݍ��{=GJ�@U�S��呤bt#-P�����5L��XTn��ʂ�#�G��OPN2�"i�(	��F9rl�-����5m�K����4�Ei����5SC�d�&(KS��X���)�4=L�Ħ���!��w-S� 8|�N> }>(~i�P7~#k��J�R���MX"&��D��ik�!���dxx�bց�8�M�QL�DkM&�$f��:�mj@D�	7��My#�Q��	4H�Vo��6��+��Z�͇B�XгX+�o �?jK%����.�[�y�k��.8��rTT4,U��Z n�����#��@ڤ�+Aؔ�a�bKqA�6�q��Б0�.i�lӋ�O{� �L5��Ju��um=<t����P~n�l�L���kp1��M�ԪՃ�'��{x����$�!��7H֌H����h��v�C���ĢQ�kR�jC+������4���!s��J�<�4`p�HM�W�r�%,֤3�n�S,����ܼ	aua�j�6�[r�1��!s���hI���¹�ZV):�F�Y�j�."Q�`�S8��º��W_
��b�OR�I��P5f�S$Q��zA�t)�wR�j�P>i�&���o@�,��w{zm<���b��&��UBx��@�h�;S��T�F��ҙY��o��M�����ږ��M7 ciCN��y+��1�w?0:(	�%�|�F������x�Ie1�'�6�G�:5��y�a$<S�\N�6�������'���$6���G	�%')�����6�L�6�v���}k�͍{���nK'u)H�ҧ75�R@�
�S�GJ�ҷ��K���mn�]F�chR�[B��+9�H�<��D�.�զ�;�&dl�i۞~��n�"�,m���'%;MԷ,�~��y'���Ph�ɹI4�ʈ�;�Gv�Z������j��@Bg�a�	$�%���w�� ڌ4��Vˑ��1�j�)�j�J��R���""q{^�"+��-R
�2bJ�*��h�BH7�v�vבM�kH�o��tѥR��L��$D�w�o]���4��#�^7k���I����5��5��D$�)��#s��4%:Z�	e~q�:��d�V4��ұS`�� � ~�v;�ަ�{��ֶăˉ�"|=MN�ӡ�5�h5�h6�h��j �ǘwa�y��$"HĐ&���N�������Ԓw @�<�4yh��<�dJ�I##��+<��Q��drY���#��vԒj @���$��7p�`j�#���ޕZ�;j6ù�$�I+JĒ�$�7mF��	�nw$��&$k�5�rI�ù$�H�dm��D#l4� Ya��I#@j�#���w�mN��#|~~D�+�ܕvD��l�[7Cd5�a�e��s��1Y$V>��Zi�F�@m��~��F#I�!�E�������6�m]��!ز|Yp[�֘�c�\�(�%/h[<�P�О�]��	��ޮ�R�΁ԧ͋��8�l�STM젍��ܸd��
aweFSҮ}@�&���5����?oI;�߈�˘;#���^DE'��]N�R��V�4�|W);��ֻ�M���^��I��`�h�ɪy��s�4�R�@��L?.e��� �$�K#i�aI��K/���|H T��!a��-}(08�z���F�z�Op�w�%X�
O$��`�Ŧ6�����k^&V4���T�\�w1�Mkj�)��ƒ�If�u�0M������[l��]�JyR$(j�O.cB�M��!�B�TS�@1�t�#�|l&&�b$ƽ��<�o[�u���PM,eR�I���,�N��`t©�g�001��oT�Р���t����y+�%��v�45|��� CR���\c:��Mh����Ӊ|��i�iu���X:��n������h��Ʀ�u7Z�?H8N����Q:�u��Z��f�x��k@�
u� ���|>w��>i�Y�j�IC�)�>K6�
vR��N���u����p�C�ahZ(�G�Fu:��B��S<R�r�%`8p�VN��x_;�r�Տ�V[��hH���n�=�q8^sr�d�udV;����+T��q��`�ɽD]���e����r�LJy�b��aC��&���P��$l��`o&�dt3Ȧ@�!/���x��VKy;)�5��d�m0>J�|�wή&$�m��t+^mP+5�dڐ�֯�	*F�_�� ��r&չI?5]��gu�r"m�`5��S��2�HQ]�8;�����4�5�Tb^�	;Q�d� 긮i_��Ѫ��l4�RD�Pג%*T`�}"oO������ޖ�H����v7H7��E�$�V:�[��POV���St	9"{�.�\���'�C�QM�:J)�_�̐����ഔBsx�Za������1#W�bQ���5'��@�4�MJ��Q�ԍ�"{�2�m9���M4�V
w�8�H�&�8�*c^:в0���F�n�CȖEԶm#D�$D:G0��'�j��k��t�b����tM=L��K����y�w�o��jF��#h1�6�In�$�e"�SZ$��պ�,MM�9�ޠ�O��'��A��s8F�6����R/�ũ��V�e��J�-�	ͫƔ�ꐁs��ڐ4^��y����7�G����N�H��<��w:M�o������5�")4�N"���B�jL>t_�X֏4D梩e��H�dISj6�ZGoH�B;|����A�ZGmD��E�"��;�U��Jk��rI�+#ebIܒڍ��^7mI'tk��Ѭ;�XwF��a�ú5�tk��Ѭ;�XwF��aܒS��-��x�#���(��� kA�:=���r�.s�Tv��GaG���f@� �Mjg����;d��N$n�i��%�;O��L~>bxġ�O~�߮g�G-�ǈ�v�9s�����A�t�GT�R�"Ge����Dj��j��rO2��q�A*�M+��#���b
��OZ�6@�b��9�9�$��5�����a9꘩0e=+B`�q�%҇��V	6Py	�Y;�6��9Ѿn����8"���\ p;�)��4HiM&�͂�i��d�����`� s�z�D�#T䉤��'��C΁59���A��P�֬��M�e�_�S��o�̛D�Ƣ@�#��i�A��h5��3�n�������ub6m:,���2��h��6 n#��j5�ۦ\�IZ%8�Q�UY��˪�U"D�1L�\eR��9[*'6��V�2��&뚝��pO� N�f��l�4�E#K^E3��i�@�e���H��> o���!ҡҢ����cTx�ۺ�@�#n/L^�Á	�=�P��x=5��8u����FQα�oLhq��қ|��� !W����n"а?Q��@M�	���_Bb��qS�~MI�'���#P1�?�z��#t����I����t��R^���������N���t�sF�x�����%�WqmՍ�x�W�E �:�d0����ө�+N�����R��;��K"X58�n�'$M����7Rܟ��Q��_<*��KC=�@��Z��i��7[s"l9�
΂E�"5�H���i��'���o&ð�%�^��y;]Dm��e�O4���w��*t9�,���"7�M��R;8���$�e��`��'�ٽ<uSZh kA�
u��К#$�5r�$�nMJPl��7p�ț�ASrLGoF�A��\�V	7��,S�	��p�m[��쬒F�͢F!!1��m;�����:h�n�R��-�0��"b�=="�X�J@�o#�@�}?i�5�K�������?S���VMRyѪ�mK�J���;rD�c���D��S�+�E���/�JUbi��pZ�ͭl�H5�d0�|�bb%�d�n�%�Y6
T<�y�l]�O�@Ѧ]iN����ZH�qA��oV�Ջ�čqd��z:�DH��mNz�$F�n� �1�{i�J�:���Gf�~dx�mo��N�blR#N��"#�!!F�j��c��x��֏4Q";7�k�L莞Lt;)
D�#�e#��B�MV(	F����#r5��Ar1�Dk�DI �i�Բjy#��B��ִ�V<ځ�:
.ٴIQ��q~'I<�����U�H�j$q4[��d���e��������@�Ѝp$�		�C������T�5��ȑ��Њt�����F��A4E:�k@ҵ�iN��
Dmb'RM��P�;5#f�lڍ�	-j6m��f�٨vj��f�٨vj��f�٨vj��f�٨vt(�Gm�Cz6п"@��ZӵT-7ڃ������=�y+�bz�7a'�Դv[��M�e�@�C�r��9����>��v���-6LY�L��߃4C"��b�[nӌ�S��6��*sP�d�y� ��|:�_��oRB�DHT������D\U�pUQz�L\�r��ND(�m��72T)�;�#���OR�U�||�>{0{{7Z�*l�7@	�*���f��I�X��w�&��K3�`5b$kk�M�4S��]��J	��eA�P(kϗ�!'��dܝ,��C͕�H�ۘ����8���wy�u$�*v(>����'�f����~�YGoD�,��Nb#QH�6֬H�K�A2�3u��d�S)�jU��!��lB��˪<z��B&%UhE\�D�ʑ.<�V�N��G��PZפ�\˰�0�S�.@�V/'&�$�3r�Q�
���Th��;eB�P'փ%�.J�l6
��	���c���׫��CW�V�C�~|�3q�L`��G[C�����C�X�!����������>|�f���Ö���������Lhq�hX���	��|+�)��50�X�Á`����*���>5:�
Èx"ԑ�1�"ԕ�;i%7�ru��8"Ԟ!�\-,�M�f�n
'���?�u*��ogZ�\�����1G Q�x�zi�֥W(�v�hۺ�uc���=�)ě�d1Cd��y)��Ѵ�_bZ$�$.��Рqq�)@?
?l(6T��[+m�Sժ�P:<��#P�i�Ls#R6H���ŽOk�%�f#w�L�~ڛ�GK���m�0���j�smW�cű3��N��2�)�ʌ>�SGv�9�S��O����e��dڤ#4^K�y<�d��L6Z�Ԓ��9�i���+�E�f�X���i"H���zU�4�mk�����Jw��ے��R_��M�10��x�ۖM�u�9\I�JF˧�^Ҩ!}�,��]3c��ޘ�R&5��ߓ�Zm�AC۠�RȶF�i㫭��±��4u�y��ƀ��l1��MfM��y!�#���&��Z֙Xt��ZOyԃ+c+fZ���;��4�EG��U#L���b�Hm55D�S��y#K�����j�.H�\�Se���Dd˝�ؒ4V.M�1 �&�ڜV+���0Dbo��h�.�!�REM����G($��QԧB�D���|�� �!	:�؈��kz�/�J�**F�#2&`���)�$��(D�"\6'F�RC��˃Q�JmY����.wp=� ˁ�]���!�R5C�g�I'�:��H$0�:q�j��0\jF�Y�Y;̦�CN�&����@�V�@�$14H��Ez���n�*h�Qdx�m�čcjD��N@�w���2�E��ВU��	"���ב ֑��#cZFƴ��x�#c^;kH��#��vԎڑ�R;jGmH��#��vԎڑ�R;ZGR΄V��q�mrH��-�
�S��Rn�DأZ�Ѣ`��;6 Oh-O2TR*z=����- 65��u�V�z>��\���w��G�Ŋ�`Sj�@Ӈ���IW.�J��%9��屳��JI�Yt7}8��*l����ש�4m촵i��t �-�G.��Y�1���]�n�����ED����&�b�Š�.`hd�O��pF���!�H�0�sa4D�$�i�Z�������*Y/Ԅ��L"7X�6H׫rb*�
I#kxSF����	�Dѳ�șr ͅ;a�q6���8������zi��ͣv�S�	���i$Ǒdt�N 55鉢��&���0Id�m$J�-�Kmi�4��q��Mo�
b{|�R7�E!�uA �M�:���� D�%J�KfЩR8ʥ�J���!Tи�Q˱*(�����VK��L"Oo��2�1G��	��s�I~]ꍔ�,����ŭױ�"&�c.r���p���Ϯg��MVʁA�P�"��LY�]Akr��-i�"m+8��4�dj���D���j"WIm!X��1F��ko�Jc��f�kJ��$֕���sxt1,�-i]$t'�@�z���o����t,��Q��NHɭ�L��o�V���'���ő�L�oM��$�k�ɣQ��m[�#ZlX��f�ҥ6�V�CSr�6�Rr��uIii-"�4�&!HM4+�!t����1�Bq�xRY�Ԅ�cjvmǚ�S�Q��˓�s�!���wmNƂ���]<_b%J��4TFU.8xb9v��y�u��[vj�������iR�"&�.RY/�-R�8I�57G����r�pĝ�"Sr�s?�����ӽ���[p�l���M�z����r1)n�4p1絑��N5F�{6�&iMG(��1�y6TƔI"�⦘f�"%��|ܕ��I M��4�ZF�NI,�X����M�D��m��7�k�ll�+|H�&��L2�kF��!5��5��D��u�f��ʊ�;�-	�ͺ�@f�{���4l�{j� j��0r@ӟ���G 5�ъu�nM��e�d|eL�j�0i�9Z�#T�b0s+	��H�;U	BY��xI�6����U�N�	�i����$�3IL��By��%!�M�%�:�7m�uMҤ��ooQ=�)�����a#j�]�b��Qi�6�C���d�v.�M'���A�f�Œ'��l�����tkS��q���uqd�zP�nݛ��АT�`�%�6U��B�4T�s$~-7TTP�~�� ~nȓ�A�t��Pۼa�@�5s|6��D��Փ��N�����Y',� ���H�S��؍p
6C΁4�&��:�o��jw�4��i�O1O�����<�}7�GO8��
(�8�C�+z�Gk^�N����:���(���w e��3�x�M��{���Dޑ.kȐkȐkȐkȐk��ב ֑��#cZFƴ��i�65�lkH�֑��"��V��בZ�+^Ekȭy���v�N�"����6�QQ���$�X�t��F~pt��98�
����%<�]+t �Ƿ�U��2ր��� �y��ˊ��T�c���d�)��^��m5��2�m�ߔ����ۂid��܀���<��j�����7 �o��PI��N@$(��br������q��s��C�'�4Oi�C A�(H�ז���6L�l���E'��2����ڡ���,J�>��A!O8��0Y��Ju�0�@tw����Rd��:��#"18F�0.DL_���x���x�4Zu�@I��Kz�����-�ni�������0X��Pnܵ��	�5F��23I��ԧNX�*kȒ���Gq���D�G+;�H��������L!)ԋ%����LcX�4�ji�072y�'�M���dR��sU�2e�
��
("b���K�J�2�T�-���������ɠl��
�N�-�->��Zu`I!&�zࣴ^ˑ���%;�c����j��s�g�����kM��b+�u���NqD��n�	7 �e))L�%��ݼ��m����E��ܴ�V���`�ó�.k)$⻬а%,�M�.k)�W�0j��OI���r�4,	JU��u��SpY��:���GgY0Г_#���ZH8N����7�Ʀ�_ƶ�"lq�m�E ��OĮ����D��x��2P~�Qڒ1GjKC�F(��H�n&��vZ�j ��&��ъ9Y"�mJ�đL�|�F�n���	��9�~�yPE23a�)W4h���t���.<������l4ӖۮNN���x��y7�F�6�xjYz���3�ZT5Y'��҉	�k�-T�C�8��R�H�5�#C&.p�5����ɣ���@��BH�ԧBG�hܘ�>*.�}o�OQ����'��ѫ|�5��ԀgDHՁH3Z$��9��"w������j�roJ��=S�TͫL��<�l�V��P�jȵ~w7vp;�n��a�4������"5P,����O%���kcSN5Xؐ֍1�S@$ 3H���]��0si��Lv�؞��X�L��kM�J"j��*H��&&�aGQ9��m����ke*�B�r)�:7Qͧ�ӑ����|���8�[T�[7I4ުF��j���rk��iz�^I����I$�騌��H�,��������EU�&����lo��	���M�M����ҝ��I-����M�a �Q�T��0�N |ؚZ֘Ԛ`HDő�ڍ8@Dx��Ь6�8K#���2��rN K-7w��H��&���b�Z%7Y���f�?�^��-�!�u���Q"-���[�;��$�[kZ��AӏRB�%��đk[R�t^u$U�$��Grh����~��p ��ש�B��N�}Y)݀��
r6�l�6&�ll�i�No�Njw  1�����x������ޝ��Q��je�a5#���I�4I�4I�4I�4I�4GA65�lk��׉��"��V��בZ�+^EkȧA9�Nt��A9�Nt���yd&�b[Y΂si�*������A�-\@�([aSd�M8���FѴe��=�S��%Ph\*�l�m��~e��F�\���d`�����Z:�"P?%�HOM�1,��;�S���a��ۢG�dI��iO�f_\�3�ǅ5J����K 0��ArO.��y�mp�"��Z
vsN{>��pS�����M�m9pg������v��rY;=LoS��4��^6�p6W���@.r#l��Bv����РL�@D�*[( ��J�:�~�>y6H�҇A1$�5���1K��i�'5jbYN"p��+M�"F�bG{�|�rI�y މ�&8 �E�Dk��5-���OS��,��#�ZmM7��Aika�Ȉ�܈�� a���Ҫ�3<��AA��ނȨ�CB�&"h\���C{~�] 1���(�M�b:#BD��ݽ�6�@	9/��&S݅#K[
w���U Pn��o��ȧ�B��'9�����	��R��Ń�$׃V�3��C��-L`�����������_�1�>k�@��8IA���|��u��'���:�#�A�?(�#��r8/������`�1�wQԐ�����%>us�qim�&��v��oA�?�iM�C�0r�"Q��0��Gm)5h��|+��pQ�O �|�W�q�lZ�\K�X+��M�C���`�m	�hnR0��"5��Mˬj�_$�M�U4mG7-�?$o��bi��֫��A�ib�_�h"�9T���+�Q4X�p1�E�+�.�9AA��l�mT��6�Ll���s8`~��_��9)�I�$�M�.F}z�_S� �:��D�Gs���$H ����`]�"{+	'�������B�J�7Tޔ
;�-��/��XZ�mN�R�e�F����"̤�H�G�rarS[;���qAId�k���P�A#��|Z$ܵ�jC�MB[���qI�[ֵ�6H�j5;�
B����j@�$�>U&��+��%�^��Gw�� ��#�5#B�$F��ͅiXɭw���7_���[M:<���d�:�ה=��ߌD�!�9ٽ׃rd�Zqj�T�Ϯgg�LD$qN��E#Ę�"�C*Y-����ִ��ž[2b-vz�6�ϓENN��6��"�UN&�Al�H�'��D��Բ0�F��7LR$�F�X4x�<|F�FD�*P�2�S�VMy���b! C�����h��S�I�l.:7��#��N�-a���<�['����cs[��.6 ��T<1�P�����Ujɰ�V�\&2��Li�`�2��q�I�t�q��Z�� \~a-jͭzbŭn���<���&��YkZ��d6@)�Dy�ֵG���v�H�`�y�΃[�y�z����&�d�T&Fx�tl��NEG��Ȑ��xgHIH�X�$_�0T��."S�_��n�ãiJ$G�A��0�$�afY0o��)
�)
�)
o�oJ�: t(����ޔ[ҋzQoJ-�E�(�����h��*�����h��*���,�����^Q6�Z��^omJ&$kCj�.�08F���9SU�q��~"R-}}-v�2��rV��>�4ҙL0s->j��P9~j�D��ow��f�H�H���J�Ci����&>��l�]�dNI��

����� >#2�ع'*At����q�R�6"{��+m (�1�Ůo���	��U9��{0}{$OP:�!&��ۣU���q^��O�����a"Ng����G��6,����ʜ��j�l,�S&�!�`��ls( �O{-~ ~el�c���=p&
&��ɯV��4�V] R�v�=�jl��C��H�kM�ȋ���^���C��4�����\Vy-���Ǩ�ud�S���{�'d7�O��8��ZnЎf�)���:&��4�TH��,b��&"\�
� �O.�] �q����$%�����H��4��ju���y�DT�Z|М�'�4��1��4�*i��Y�ZZ\ Ni��	����{L��q��#jhu#	(>H$�w���и������!V�8�Ts�F���uFQ��Z�L"u��VҐ����|O���S�m`uF���`��Z�M\�V��_��S���ɸ�BǦ48���Q�p�(�+@�I�C��S�� ���u7b1髟�H�R."�1����NS?ɍ��J�1�.����n%v��KS$��c�~փJ�&���H5)Jd�{ZVnN�	!$��4M�gѲ3�#�yUR�$J��P�a��ؕQp��m������U� $��8�S!�����4`�oO�����R"�$�6O y4���J�p7*uC�|y)ɂN�ih�43u���b�4��$J�,z�U;����Mi�x��"OX�Z�b �#�K!0�ή����SɺRo^��간`lmM�M�i5$��n�Z(Pq1~��N<P�`�0.䨈��޻�ޥ���6�<׉8LRBk��ֱ{S;��%g�h�b�1Q�����T�H7��ƽޯ� k�)h�֍�(y�e�~�i 2V�.�������ja)<�9 �rm��Y����Q���<��)>���։����:5RGeq�b���k�ã�=���5>��M6�xL��rF��>ww�)M/��4S����5>��������ڻ��ĒԬH5w�Ǔ�(.8�i�{I7��C`
�_�I$�i#���B���j�l#t=����ǎ,�������Ԩ�"�rH��Vn�3C����lݡ�9B�:��M�i��.Jg�a�����-�=Z�g�1 Y0�H�t�H� ���6������"�0�&Vk��ʗ4=�.eH.N�7�I��Ʀ��D�j��e�$wz��3�b�i��֩4�W��H�()֙�����1�03���-��#Ku$#Y9��A����M"#��CC|`Ēe�*D�*D�(D�(D�(A�(A�*A�*A�(����ޔ[ҋzQoJ-�E�-�Ŷ������|[o�m��٬O��Rx��sh��:��H��6ydZ���s���5��1��[Tnn�T�?\䁸ځh�sC���,/sPl�$z��30���*��>t&&��Phca-�Jn��Z��*��oI�sh�Z$��j�n�l *#{*�i��
[��4
�shc������=������r��¯�g�ӌ��~n�l	&(8\�E%!�h��lk�	k)S��r~q�l�{����S�0Q���(�m�lH��n��^�7�#L1��j�l*G{{}.��z�|�p�d��O&�\ͤnF�kS�"2՛��$�"%����i��b�o]�ͨ�9��T��-��5����̍�'8C`oQ%G�t�U4 =��. 2�Ԫ�c��A:��%=e�Q.Ar�H*ET����@0�*P�.@�� h�h��z�A4��-7�/8x3e���8����Oh~�|݌2�I:eE@�ݓ��;<�~:N	-J�$a]"JnZ@(�$�&�&��"�Z�Ƥ%^Y5���!	L�	6�B��kH(慁(�hp��	�ޚT��nڒ�ő�ֲ;��%%	L�!)�����I��������$��9d���J"��Y'7�#���WA��	D�:ʆ�R03H�W+�� ���)��қ��Bu6�ā���!,уR�L������]&V4+ Ԃhj� kDV�S��N&ژ�*O[�\|�_��*>(k��s�4*� �rꨥ��#� D�pc��zcu�|nT�(?i�{5�A��!k|5YI$�iIj֖I�!�i�ɷY:k��n���Au��X�$M1�n���I��	�4&H�lI�l�"s1��s�"��=��7hp6GJ���A�| ����"5���Mgs�j�֒H����1@i����	;H���㭇AfS16�t��u�:$׻�F�#���$p� ,T+��'�8�`t[;�����e��I��"�o!����mn��c����i�iːp&J����9,Hb���4���Z�O$��jG�ڲ5Sz��NDzӹ�SBk�T�,�1�ڨ�ff����>l���燓 	�ln��&����.	���R��E���m�m�7v&�<�����n�j�#�Pcڃ��dŨ׵9Ш$�7_�ed�m���0��l��$id�:|<]�ڶT����Ϭ"T�Dqɪ�=���T�`ݠ�'Պqi-��~�C�8xL��x3t�s�
����e��56���6$�e�i�I<uQ�A���(h$(TTT�����w�Pz�$eq"��8��y7Z״�ٹU92�-T�kϊ���E�bO��m� ߋ\m��`3*��5�	#SND
pM����:y~Z��l�I2<�mGR��F��V�*bĩ�s{|akH�,��
�±0�L+
�±0�jBڐ��-�jBڐ��[�zZƼ�Щ�kF���$ot �*h$LD&�@l����a��
��8��8�����Bf���ˎ#�9�@����%��r*�+��Z)�ij�4�7L�7��E�w&�Cm8iő٬���J|���5]�3�P�z||<�H1�$��n�^�@�Tisk��i�04ø�A��u2y<�c����lT������6�{$P@�4L2Kh$�i[��3��H����lѣ��� w-;,�'�$l�I�f�#U�uH@��v7y5Z�+�94F��*�
���,K[nt���N`2�}X�=�ȏ6��Ղ��z�:0:(9�	=\����F�$Ѻ�����Ue$�i6���7�sj�u=Sʗ!��a��d���|S�x����y��J�hEhbbQ.��CD���'�=����%j�TO#�Z��[R8��;>��K�{�D�Sa��vO[J�1s.M�ɂ5��<dP�v%T)m�)��áMfj!$
�P���F�N��	DK�M˭L��� )� ��- ���u�D.۾	�g�܄�6��CQIDt�[�J�$ک�������y5�u���ړ�1 WH���R�\u+��M\�zi�SZ�[�L��^qq�C��E~�x�2P~���h�т%����7�L~H<E����5����x�֡�Z�I�m��n]J:�8V�ϒ������vH�����=@a����y�&ĉf����]-
��BCCй�b籉A{[rn�S�H�)�ݕȑJ���P$M5ZӲ�Hܦ�	�i�����ĊЮZ�rL>T6P�&���i I$�	������u�m��lH��� :��E`3`\�b,�����@ީ��D���č2֕&V(�I��u�xL��J�i�I�2����w*;�O͓��Q1D�kU��j�����Mvz�[*E����x��v(N?l7����u����b"r%��-�ռ%�d|p��M"�n�曉N�RFȚ#�ˉ�
��;�f
cln�A��6`۶���Y-L_6���9m+|���X��}?�;,[h��޶/QQ�Oj$�p9X�
l6�C��w9�{d3z�@u@��w�BD� HkX�T�╄���d�)f޶A�V��I96-j5�V�l��<Zy����#~N><P<�$�L#S���s�1��Sa�ۺT��rid�l�S�B$琠�p�D���[Ƞ�:�R'� ~.�D�T\�ɽY�VJ&�b�D�9�>\ף@)�O#O�00cLoL0�� �z��@�$���L��I[�Bj��PJr ��Dv��
t�:ې����z�Y�G�EM�zT�z�H�{U ����̵qC�ɺ@)<��B#���@xjT"F���Iũ���gx�&�4��*D$ةw �7���B%K5΂����(A�}[�L+
�ޱ0�M�
�ޱ0��-��-��-��-�
�M[�{zT��Dв"<�7D�lѧˆʌ��8�΀4���$t�Ie��ȓ�7R����	L��3Gs9U����.��x*8�pb��Q����S�4��S����k�A*���6���S�����CV$ש=D5_�KS�����Q��%�H�'��No3��#NJ�}Ae��PG<�]s�[�����"j�P�iz5��8�H&e�#�
��� \�["Y���(	�~-rkI��Hڧ}n�9�]�>�I;8�6J�ԋ��'Y?,�΄���bPМ�q�1��+3Oy6M�cɁq�D�ֆ�����+�[ѩ!�T��9��Z�(�72�78�#B%�	C^V,����(��'�.T��M����4��p��Ւɲ=.z�]�bQ.��CD���'�=��8�9���r}Dn������t
""A�m�m�M�ye�2\�'״���g`IE#�;>��a��.����vP-S���p!��H��uq��|��P|�$ۋ�r-qq&?-W�2A�u���8�u���8pQ#�I�F$7L�S$p�n�4�W�r��RQ6�ā��I�m#�q^>���v�Jjag�h< �@;pm#��!�a0(�#n�Uhc>O (�C:�o�\��z�"۫���G-I&9@��H�V���f�mWX��QI�S�Z�������Q���i��C�u3ԄOk�k�ئi�5��$h=I�3u#�0�
㇘���4Q��$s��y���Am��l&�&.Dz�v�Nri��r 6WY95�f�yC|IK6��@F��F�v��瑠�6Te�F�VM�M�SH��$����dZ�Y����ji�)�ͩ�C^�!$�e%��]РOS�
I'&�y�~~	$~p<2h��<��kF�6������dt`��u1�H�58�Go��&܄�	��%!��j:�ě�ג`�� %��5���0_�Mi�$�"��h i!C��a��T�~���k��c���hY?
�=S��tkT��s;)��Ө�F�Y����ƷC�<z�~t-�y���R�;F������HTL�� ���8�n�e#�{���N���*Cy�6�����'�c�'VJ
����@�H|S_���oo���O�� �	���п�r;:�4��wv�O7�fW���$�'�f��8:�X�����qi=��S)��7X�M�S��9�p&;݊�L��Ȁ]�� ��@�bDis�y�V@T�ޙS��(<�oZn��1�Dx��P虑ѷ����ƣq6��9�����ژ��2~FƩ���s?a�)RI98y�؀P!$u��aE��R�;�5Z��L�1�PG J���D�! �4ȑj�A@�f�*\ޒF���jDjSS���T��N�-c^�8t"hX��&��U�zŪŉ�b�b�ޤ7AH`�!�
C)�R1Hn����h���ާ?�tF�����FD�(�4����072�n�'>���ߣe�g�H���
s�M3��U��{sJ�oQ����TRX���'q��n��A+�e9��]9~[O/h(r-4��4��Nȑӏ?6"��T�Ԅ�6���������jvȤh��VP^T�e~� �j�EH6'�&#�@ ��� �)��^�C1�A9�՟�h# �>�^�崮���Cᎅ
�[sz�'�S����GsQY�vl;(('�=��]��i�]��tk��vNN2���L`�f��eءٰ:�~�L}z�6�L�C��UNw�k�(��ӣ�������&�A騬�u���SĦ'�.�ETqur�C4۠ʃ��7"TF$b1/�%���(R�AV"���uZ&ZL�T�S�#����x���������ܵ9@S��;�$4W"h.pࡎ��oi�g�cB���\Ў�]���	@�4K6(�+��~�zk5sqH���s�?H��B��c�U���Z8����?�b⵴�ۀt"c��S�
?�*1��n7SSp�Z��
�7��������Ғ�Z"5�K���Q� V��Q�e�S	�N��������me�S	�`�hW�Я�*8px(�2Lr8(��xqm+�8< ��Ѹ��w�!Qޘ��u�d6��x�ͺ�c����W�1� ��/8���q%�A�	f�"zͯX+ՂA4kqJ� ćJe���P�)��W<�+�"�EsF�>���D�����3M�m���FW9E@@��M�ޕ)���C�v���M��L�>�J�o�BoĆN���4|6�~I9�N�Jt�Tty��el4�I�Z:�|D$`6�7R���)-$�;��ԏd�#'r'Ѩ�@]4Fo\�Q�M��Bc���Y8ޒH�ߛ⥳��L�#�e�F���%�@$�!�"&�=�8&��PkI����'�rjI��l�Y5^J�]bZ����	����HN�~���\���Ʉ�5D��4|m�ɭ"L4�9��U��;|�_���V�p615f��#���5F���GE]�2��#kVn���ɡ4�R2b-�
TF��ו���5�<��P�[E?h�����R�J.�X�S"JL$L5�W�Ri�wM,���I�$�77F��J�9	��/k$�֑ImV������ڨ %�*I�M����^�	�OO;������\V>7H�GB�J5��6�w;U��.HT1�T]$T1�nx��q�U���y����xS|&�گӏ�Z��cŒ֘e������!�u�4��-,�-����*�''"ց1���<ڧNz�4;�.ىDȌEO�o�k�浺	����}i�\��N�o �˜$h�GF���4i�;��x���U��A�֫��2%Gv�<�ַ[T����#f�0�J$�ؒ7bŪŋU��-V,Z�X�X�j�b�bŪŋU��-V,Z�X�X�7�
,L)#����� #���A@eʣ�o��֪}1�P�\P؎�ǜ�
�9>�G���~�Dށ�VI&��$OkK��g0���d�Uًfc0�j�-s#5=[.NK�q��%�!B��'%F�98�2B'����6��r�&�� ���f45A5T��zV�Ƅ�K�� ��l�c�7a6�c(���&�Z�@���7<�Nw����Q 'Ce�I9lI@󒪪S5����M/�[�Ki���oh���ۣ	iJ�P�$�+'�σ&9A ��]l�<I�:�ǩ���P�R���A��{b�l��4���Fܜ����\�o�\m	0+��׷�oWCLܩ�9�Q�P��i�\����O��H�"4�zP�y}hbR�*h�TK���ZL�T�㓱����Ko�EO�b`_��r2)��K�2]���E�ߑ�� y��b��y�'CzM6��%&��hQ<�'���p��5sqH<��~	,�"#����y���H<�ŨEē:�'��KQ����̔K+��%p5���
��QƤ��d��1����L��V�[q�,��1�ĵ3Ėv��N�QID5;:��ǉ�$�&)�S���W,LK7{zOR[s��"�:�F�ZNQBNi��5+�MD%s|SX8Ja��.ד�ŉ�f�mM�S�H��Mo�D�h]���ۥ�D�܈`�涔�M�B'	��,2��p���u��'΀6ˀ��{�C`��ۘa2������ �^��Z�t%���i ��ݭaP�{e��On�RD��)�DI"��t���L`�#ۼ� �c⡉�+�1����lu~�$S�M��9i#M@�̩$F<NY4�n��hS���Nwē���b[�y\LhM9�^I��n�ڽPn���HһZ�K_��6��$ޞX�H�\g�v�QE@���k����q �u<�A<�$����׵�8���	�Lry�T�� ���o����HIm�vX�_�꫶��*�5"ro�HN�v{%���b�ct0o��Xݧ�WEmTQ��&�L�H�	8cWb���ݡm�*p�-�Пk��N��K&�\�$������&��[و��,lɨ���pٖ��˚u�S�G��z{�b�;A��zz��~��pM-��BxQ0M��}7��^����dHc�N�H��&�OQ,�O�J�-���P��`d�i$v*L<�*Gj�?T��S�5�j�4�"$.~ݖ�%F�0Oɍ��M�n��
���·2�Z4x��7,�9�/ܝ
C���"�ۭ�;��p�p���a��KL�g���H�D�"{Md��k[�� K�����;7�m��u�L#>h$2~ݷS"dI['Ң���,t�O_��D�3�5����cS�HM(�u�ո�V�j�[��p5n��ո�V�j�[��p5n�$ap�EH:��7D��w�VMV��A��Wg8'��u�����Mj}��j�@Ϙ�?`�b��vsh2���*W��� ��.d	�㓛�D�{��6�K�
\�����	�U7Q�l�cM�MQ��A4�By��A=0�a�15�A1�o[ѳ���H?.�mP"�f��7��z��������# ��Ċ�ʛ�G�4ߐi��(��-~y(Oзth��`@Ib|Y ~#r8�|�i����_\����ʞC��e���S
��6A'7H����4JY{X�O��hבj�����bi��"�����_�� PrkD�%�ɱ~�u����(F�&�"OX��G@�e�5M�c�\��"-l?>�6ۨ���į��ăkbBNĄ[O[F�?�O4ZO!CCE��V�C\�B��������4vhvrGl����Oi����)�� �����ߏ
.�\�qC �:S/�F#�0��a��H��$k�ț֙!�<M�}?S�����I�6��r590��d~:ti�7�f�5�9�1N�n����oRkT��$�	5�ԃ��S;�f�I�و�jD�%����Ǎ%"qC���$;�HDN�5$B0z�Q�ޠ��"k�Z��ܬ�.&�j���	ũ�Q	\b��f�a	f�6�Y�Y��r��RHJIԑ9�m;����Ƽ�)�!��D6Ln[yY�b)#DF�	%!��ڿ&�Jt��ĩR���Uc*�
?l�-l�j������Щ�T��]����U>_���v��ޘ�?.�y���D����G%�X��F I��1G�K���=��l��i�o��Ҳ�.R4�ޣ���4�I�:�>6��DN��F�m7��@��6�ym<D�l��LX�I VI��aR5c��cIq#�B�j�C��"O<�*��M�?<���iA܀�d`�w�[nj
?\�������J&�[&���|���''<J�a�.Im[��&��L~oO鋃���I%��p󕲄��n��b �K	Z���A�p�S��K&�t�t^aj�H�����{�{r�l6�!CR9 ÊF�~�nzm7@�7M7d�l�Tq�k�$��p6����O\Ww�� D��Ș%:��b4�eMR ��!M2 �	���j�hM9!�,���ݓO����A��n�S0s�H�;<檈�hLGH<�Dߎ����� 6��ȞȞ�11�7B���1�l���npL�q!Atґ�M)�I�ֽ�>_�S��ߓ��Z��a�y̘&��\%�a���4��$�'ht�&�nn�ސ9��� ��I�mD�LEH��=_���c���x�4��Ov_�?k�/�G"� I�V�d�&�V??4���6�����q7�둺�� ����'��d�����<���'�! ��u�4c��V�j�[��p5n��պ�����>������>�O��H��݃ɗ������4|V1������7Q<��%l�oH�R��h�a�I��Txݺ����.��\�-vѴh���bmZ�VѲ(1�%c��L�?;"i�_g��ʅ9�@��f����t�ka���Z�	Ӕ�ǋ���1(eK� �|�Z�":(#[ ��mǗ\��8�<bp	� ��"lj�h0��7�O\H��4�H�H����'4&
�ܚog��FU�h�51��>k\KS=�}n��ѭ�&��dDeH|1N~Y;Q�"% ��4�DYI4�Bm7��U4@Fit(GS�``�F��-�Bw��*��ysr�X4��c
!�]��?[P0L((D��t���Tn��Z�_�D�Iݦ�w�7?�~["c�*����k�U���2Щ��0aw'#���>�����]=�q�8��'յG�.J)c���<\a���>�Ns[svrr[l�M	���o$$���Wx���SzKHI�"��)�&ł0�Q��6���U�ǦWZ�N�UJ�:�i�V7r�;-Tu�_��
�`�1��2Q8�%��R{�.�%��q[t���p�ͺLY�u��qo��j�����h����@�Z����Ԯ��k|/ͭɡj'�^p��"qB�Q�9Lb���r���<�"��bx���hogd��X>�#�5L�5�	�*�J�L1ݛӸ���9�o@ɤ҄��ļ���c*�(!c'�^̠�~��ߘ�Pӗ]2���ƪqS^�y���bM� H-�;���	�@���	�T�o�c�c�D�� ���i�|mM7��QAk�s�{U���m0�l�N|~�>hi�S���2Zi�M����2D�	�$��ۦ��&��I��6�9�T�	r׸���ؐ-ڥ����]�%�zh��Im���4������Z�:�DmS���̀҂�JD�:�)"�4LF��K�D��a��q���]{�E�6�L���d�j&�2ַV�&���mr�� ol�ؼ�Ӎ$suQ�� k�D�\�Q0hh4����d�kBI�@kk[�C�NT�)$�Ew��BP� ��q� 0��x8Z�H�Z�oS����I��%�4Ή��%�"4���7F�7�Uhb5�U�+�:�h��[3��ڔJSl�	�&;��V���j��@�-�'���I\+����$D�W�j:�1~�>Py7L�U?@6?"~w�O���	�(LD&�@L�4���H�ڒ�RE2�#��HIxtN!6JES�@�%k�M����$%���S�4�Atk�$n�m�F�D���8�F���G�ϥE"B�ɺ�I�A����voS݌G��U�٬H`���L�0R(=\ǓG�{T�ж�mM�Ქ��̠lR�$�I	>�� n�#i�E�G�8�p �>A�|������t��~�A��t��~��� 0�J��7�Ǐ��<�&�,^Kg���!��꧓t�Iȩ�꜍��2�<�Gri��З�������
]CB�PoJ�Ĩh�b�*� 2�P���� ud�Pr����[L8��NI944"[��V����evq���+� Z�"G#[2F�@��<�p����Ǐ .������� ������M�K#rmL�;#P.q@Q�P�TS������� l�[���z��\�H�l�����\����$x���4�>��dƼ���NI�8
�@h�V�|�&)j��֦!�h�9d�A�rC_#JgB#���V:-��Oe�����**?$}-0k��<D&mo�H�(9��ߛ)럆Y�\��5J�OQk�Z�s-
�q+���x�:r���ʀ9sO.��p0+CD��NonNe�~.e�����vsl��'-��srn��[�h\�OH��H;/�kn9'6�jE�&��mx�`"S8MkW�r�V�]O:�h��kG��I�n�i%51D��Aq�V7R0?I������X/�scx��!�ܤA]"Y���H�zn'���M��S/�u+��Q��n����n$'�KY��I)= �M!Ԧ_�86(���&8���֬jk5sqX$���Lm��Z�D��"SzMH�n�ē@�k��i'� �`�h�d�~�mHDd�X�]�i�B���$�P��$�4��W��4!�hJ���%.�y`�ːa5G��9��.����t��צSDdƼ��v- :�L0rk�Ry	�mZ��1%�����C�k�
9 s( &6�z���4��`��dm2"���^6F�?v#{i�.Im���i�����!J�l m-OH���u �#T0�a)h#��#Ԝtvz�
n����F��Ss�g��"���p4�&��	�`�o�&���R��X��,��591� &�Fn�k��e:��mM0"S6���`�54H����H#^ݒI��FQ��/xjn�1SvK)�������NkTԖ't}kJ����@nM��)��cj&n�mO���|S�m"X��1K����1Y$����V�!��ܽ[K����:0���ѡ�D�O�\D�PZ�ӄK�.�$��U�L'�C��,y=~�~�L+ d��T�Z1�TkN7\N0n���sj�O l�]kCJz14yX1��MI�ʕ�u:�S�ƮI�s�����<~�����t����7J�(Gj�(S�v������<�ނNY4�[���I��L���Z��VʘDD�6`��$Gp_��_�4S�5J���m:�^���vNy>�Jp���Ǩ�᩼�ؖZdI��T�l	���Ԓr��<�'���wځkAB5t���bD�A�F)�F�6�A�~������$�ؒ?b�1�#�$���L�O�S����L��.��2<Ս�`m[�޿jާ�kfPؒ.o����4v봡>�*�?h-*8|�"O��(��H���9����.���h�Éh�(� ����'�2�t&�^DG�̧�'>�����-v.�T`ЁQ�I��ӏ� 7S��*G�ӈ�K�8�Pإ�6^�'Av��EA���:e
,�&-ߗK��|�xy�ˁn$��_��ĲH��^��dm4�#�&���-σ;ީ�U#�ym�A~9vJx�Μ��N������(�&�i�+T�kt��� �0�F%t&4/��V��&$��iI�Tj$�%l,D�)�r9p�7�"%���x�8��8���B��v7-�~Gj�����&'�l��Q�ʅ<(�2�h�ڭv����L8��9�� 	����8�e�8��{�bR�%8��i�4��{}}�)�	٪���NO��@o#B��u[к���F�͠���*��p�f ���MH���вlQ8[Cqz`���p���-��x��d��&�����p�$��EJ�jk7SSV<��h.(��Mj�R��V7���$��D�|�(�4����|?�׆9���N�&Х_�ʹ���c�b�hhH���������?�-IX��O~�?ޚ�xc��M�L�n	��i'��uጥI�6���'�cV�֎D�l7�0Nj4�X����n�$4,�R��Q��\{cB��R��\��K�'=�6^���R{��QBz�t�$��{��&)d����k�§A�m�5�����)���(�l�T���ʃLe�S���Z�F��F�#)���BeI#�A�K#�S�3AYb�nSJ#����.��9j��Ly"l
��*m^Dd��S�z�t����*�L{:"Y%+#D��w�X�Ƽ�M�SO6&�T���b�)���kACd��m�;yK\��&v	�-�M	��B=�*�16N�S��E@�'�Ɣk`��Zr��o#qȈ�������ו'GS�ֆ�0ju$N�6�޶c�˄����V�v?$v�oy�&��N����ji�)�1�ktL�mӂ!yѺ��6��4Ҧ��eb���sJ@��$�n��D�ܻU~�iF�Ĕ�"Б$��0$76����ڲC&N��-�z�����T
b(�@,M3�������:�@���S�N�R�"ڑ�����f��£�e
O�*-*T�p_��7��Ԁ�h��f�oK'� gO�Z�&S?X�V�UF�A��[��mS�M-��
�w�=�9�*��N$%�6[�q���*<�6��Z��&���y?9�[.K%��Z�#)�7VIǛ����ƽ�7k�M5����F\y�ЍL������z�n��$٬���b��&����n�m��#�����rh��v�?�1�|�������NF؍�� 0T�>@��P�[���#?D�N��X�F��S8ݍI�֛U�gh�q11=���Z&l˜�Ap"��C�ӊ��jcC�áH�i6��"h�1s��[D�bj�?"}hT������3CC��6�~����6�� s3U����\f_R�\\�*"뒂.�">���i�������D��S<�����4�V���u9HT��*8�r��roJ)��[T2;ȴ�"e�e��9R{C"h n�N��gB��eMW1Bm���Se��a7�OpV-�hy���	=HMꦨbӠ؉|ܘ�e!D�&�D ���a �;M��FI.(��I�ܴce������7t�?i��J1��s44H0�ER��m��rLb�T��
�y��*�B�ύʞ���&#�N~[l0Ȧ�T�R;�BT�	��/��-0Ϯ�����t�9==9�`P@ךBM˩�ڕ��a��1������U�&��R�I�0wf��}k�ƱhhC@�
�_'��郄_9)�>O�����6�8��:�
�н�joB0
�TN�X�zkE9ja5k��^;Ru�:�X�
#� ��N��f�n����V6�*A��w�ͼnP���MH
�h��oI�ҲԬRu�J�q1�Y)�[�չYT�CSr�k��
@j��ۤ�&�6��mA���HubY(t5�#H^]:��Y�vɴ�dy��֘�m7b1�"�I�TW�A�R=������eA� IR�=�6Mͯ&�YH�~Z����VS��dӡ���nߥ�s��a��&�T�ճ�=�7S�4���H�����2��	[&��T�ʖDN�4��t�@1��zT�Y o���B�aY�iS�S�T�"C�ii�N�:�;��!�!Y�"���F��4�ҿ:�G�n�"(}�]�BN��ގ�eOfI�v�HN-H��J�'�5�~j��ĕ ��4�ؠ��74)/$�t><
�N�b�����;�AQ9��B��A�z}�(D�6�����%i�1��0��a ~ht-�[�!�Ę�&����Ic�$O�{���"����m
�BR��Cr�JlyM��F�U:��S�bا<DNrY��h��&H�=�N*~sl*[?<�F($�S�	���8�"�B�2�v2�L�탡h�u1j�0���̮�L!�S���V��d�%n�C)�����M2aӡk��:j-sw���Z��^�6:5X�Ӎ�4�H���a�3��v; H�'�Jdm���蜱5��(��U��j�17h�A�&�Ȕ�8`�r<�[.�[sI6
v�{�A��3A��E��8P��F(��?7M����&�,�޵o���3ijc^�|�s"o��M���jF�p9/ޯbDfGZ�	�bm�52$�D~�������2�Lc||��7T��'J���i�.�Nٸ ��;��i�;��y"_��"i��16��nn�7N�S�虂St���Ʌǚ���S��sh@&��N���QUiZ6ZQg�S)��e��e�"�f�k|H<ސ(#[��W�C�櫼�StC��@r.������pe�܋�33@�p��6�q��p�N\�"/T��ͦ�]�P�>�.��g��1�m������d�Ջ��r.w7r+��먜�Y��	9ڧ�=V�,S���W��eꔁ�i���A\�	)��#�Ԣi���F���Ȕ�P͇4v˲�;�
��s��9|em�ZVi�܄�x�^p��7�6�c�9L$KR6�z:ۘ�d�N�F���"���ƪ'g8 �Ϝ�D�>����er9�NO�����$:���UV.B��� ��H�*a�E�˗h{} �Lsj� l�
rOGsN��?"F��'{{2�	rs����bI$D�_�Ϗܝ��<e�0M�;��ƇQC|5I���2�HNm��В��v6��&�cx6�'>�W��J�i&!��+)Z�ɭ�4���Z�kZ�d�B��vq<�u�D$�%��ӹ9�i!/��������q�]`4)HcPk��hx�A���xS��at�d��6�ZF�����2hI�5�SE����4)�5�Y%����"�Y�!5�ܜWu��j�HI±4���A$i5�ĵ*�\C'������T���e�Q���d�ר��E+x6R'�8��t���(W#��\����"�c�hz9�.a�mQ5��P�u�ar@I1��$>m]�'Ce�|��-S�).�^6<�-y	
"a��ni#�"s���<`0�M�<�3d�0d�������e�M�01�<�LR��"aI�CX���$�l1�3t�#��ؘ�M�k�r�i��F���ʑ�RN:#S�E�U̍�d��
14PP�)N�Q�l���`�'6R�8L�޶Z�!�ܬF�&�[�����S6�$�H�����B��Ά�r�NS)^����G���)�����{9�Z�A"I'M'�+D�l�U1BI��ܩ�H�'#j0D׺ɨ,S��i!&�� M���.@m��x%�LᤡٷR	�HR�4ɡ�,�^O�b'{�,zZ��[}Y�Q����u���cj&���m��P7~l�4??T(y��(�@��Nr)�T��;`���\n1m��~w�\�%����:6-h�R�3H�DL#2ڕ-�� ��' ]nm��g���8� :ly����SG��B{jiz��&Z�25�x��;���~w���PTi�6���#R�f�˔& w��ZJ�e:{�����m~��@�T�'2�"`���D�[j��n�?����H�&5(w���s��L�16�#5L�;�IӹS�b�:6�T`�P��5���2̍�#lȚq֝�F�D��j�z�*>@u�F�G��V�y��#e�M��~�z� m�ۨ�XD�`�e�m9CN`�?N��EGm����6�S�����H�k�����;9 qR�Z*�\���)�e.OǞ��F9#��۴��Eݏݏ���M����Uͪ�6~��Uc�&��b�R�w"�h{h�)��^�4�ۥM������ʫ�c��tS�J���(iPJ쎠:~y1����Oo��@�9"p6)���i��CbT(���i8�lȅT7,m�=�F������DH���FA�) ˘-�˥"N6��Z@mX��Q���Q� sL5�[��@�y����bM`��Ef��B1&��CR\$F�z����Q�=@ ��@����|�t*i�j�K�T-P�.��J��e�R�AK�AR*�k�� ��H�*a�E���4F�n�l7fF9�����6�m�wg����:��d�7I:�.wx���z��`u�1)	f���4֤+��U3��	+�PjL�y�/�iD�D`|vH57����՚��Q��Ө&�mBL��/!e��,�ZJ���V��c�F^B���q8C��)��B�L�?���B����P���$]o�&C�Tq�Z�ZG���ZJ�ҵ��U�R�i1�b�����:�M�0�BH,LK6�����&��֠RZ�hVS<[Rz��hV)]gP�`�T	�D��&����X��F�R��6"'�	�`�č�f����&�ːҞE]DSu@�aŷ�9�O�-�8�r3L{��H��#T7�l����W��̻�DD�m��'$kպy͉S�8�I#$@��H�H�j�l���	�6]����/S�"����Oy��kn�R6V5��D�9aBbs|�<&}KF�(I�;�;
v"?}$l�?��d�
��VR[������Z��,�H�����"� \<�i�_��&��k���BiNɦ��.��܊k��ؚ�<ڎ��^�����Z�N��Y�o�W�Ϸ�P[t��J��e���*v~�ˡ@1H�9w�"5�DOZ4��k�I�j���!%��� ���QC�0M�;�T����C�]�~�:)�bg+��M�V�?[Y����bT��9xb�'F��\N}kH��	��&���w'��aRڃ%v)������M��X��$�2��0�:�K�p���;_;����kV�D�08&�����a��C�@���#�A��&&�m�"y�������f:�rP"2����n:֟����-�0ū�� ůPɍ�Sn�~X��Lhn���~x���5({;�F$���#��N�_��@����7KK��Pi�?$~���lQ�.�Ґ��.<�)	6�!%!ܠu��T$�n6(�L�d�q�b��#M��������#J	��*>akb`�?\~�����7`m����$	��MS�����hǑ����k��1qbgꇚ��������vO�'ۭ��4�'�6>Gl�7g��f
�@2͙Ɖ�֍u��WR�8�|����]t2s�xyN6��{���#�P�M�FTT��#�<�<�x���QNe��b�˴
D\S�NQ��Z5W&����0n�3�z�[ 7A�AH:�m�mj��Q�J�5��f$k�Сqqw�`��%��Z�?!:;ӎ=S��'S�\� LrS���&(;���h���*>{}z�J��{����U�Q[T��ժ$�mA�*�k��B5�H�,�Ƥk�E���iN���k΄�A�Hb+$��Zm���bm��Djkkn�deEK ꅡrTƅ�J�������0`�"��V��r*D�R�hD\�ɚT�q�\��6S��Z�772�������vPOO(*0R)5Z�dU���ެO��@1	�X-T���M�)��r�G)������mM�i��H����p	$[�	��+��ּI�V��I�)2PЮ|�2R�����P��"V>e;RV>d�:���ħ��<Tq�"m���
<Tq�|����S�Le2��^�n�|�5�kp��a�-Lb�]hi6��$�Įޒ׊ep�NY��ķ�ĤP�'��f���+��(�4NQ��0k�hq#@ժPG��w�|��C�H��"D�-��N�&��y���`Qb�P.y����Th�ӝ�O�&V�Pd��v��T��G�5\�9?=M�]堈
�CdjA��5m=�(��z�4��ճ��0��D��8�"��|lM
"G<�`�?F���"�A�~6b_�"vNp��qQMN�t$O7���H�j� 3��H�6�����(l��ɥ��O��=��,�\�S��ci�m��M~�Nw��f[��h� WkҤ�)Ǡ�HDTk^�n�z&)�il�������<��5p��ԒD*�;�G�VJ2h�6�A��U�U<�ٗ�Be4�i����EF@�[��IbD�58����������r!��ߟT���\0]���h:ѡ�������)��ҥJv�����ZP�S�C�2L�	J��zŲPkk��bKgA1Do���҃�EKj��nE�\�&��q��t� k�زF�Р@"S�*~h>.�)�0��%�d�M�i�r����4~	d� �OA��s���	�����it/� k����ء�n�M%��F蒹���Ū�M�#Q,��5�Mk6�jVF�,����c�{n�0H�
���l �0Z�������+���Ċ������ ��T��\�>8�n�6���h�-�&1A��	�	�I���l���,V�	�J�~>c�Ur�Uq�%�)��۬(i�:� O`�|���-LD&T����i�����(r�;M�KV䉋���� n�z��p#�AIN�Oi#$�EI҅'D�䉋�[����T�
W�q���U(ghǻ��t��$r׸f^�-��?GD�E�h *����S˕J������A΅P�HB�Ў�)�b�WF-��(��c�crtt�y�sUɲP�T����J�?.h��������)p�V\昞��sO7l��±��t�d�6����0;�	��a����ԭ��U#( �֏A�E5�x�&�N�C�Z��m"?kH�)&�V�v>�`��"rX��7r\�(1���_��ڦ׭8�=��m�''z���P�Uj��
my�P$:$�_�^��Q2�4F������x�m��5��$6K+'$�菛�c��s��SJ��Y�@��K����\�t"��V��r*D�R�h8 2�ʀ T	킃Q߆;-��>�l��m6�e�	mɰZZn�p\��l6.�qG	�����^��:�J�2��S�d��h�!&�"lQ(�f��+�@��P��<^�A�֍�F���~
�Èx�� ���:����η�Zu= (Y�� �~�η�"c��ML���S�9n!WXDJ1�Ð�B9ň��%��_��1�^�:�n���V6��%��oI�'���i'�V�i`�n&�Q�kQ�UᎥ_��SS:����?��hu�8�F<���DC>#pfa�+����I$��ΥsUf� u:�O;�@�nD�&�s歡���-"\�hNG8�qU*Ӂ(&6ڢ���02�Cgϣ��ci����U�D�P"n���@7{u$�-:5���C��#}"y�в;7�e2Ҳ5��n� PM6�&`�DZ�ڏ)�Ƣ�����S�u�t����J�<��'���5�#)���E������z�LI=_H�F��"�nBF�@�9�L|m$;6�B+|�ejt(n+ #�#Q%���(F���Z�b��|� ��l����aJw$�9oQ�CU�zh��5t;@���^NJe"y]N�w��*�8�f�4P�M6�ő�!'�cI@c������6&y�%�N�D�y수�-M r<ޘH�kȯT�>+i�H ���0&<���#pMx�Ƽ� ���mS�$�t`֧r�Y7h�S�	� �E���H��:Bne�Ȝ�h#��O����WB��(Ǫڜ�t2T)8A�i�SJ��N��[���ꢹf�@��ĪYz	�
*Gl�����oV���ו#[����':	d�OW�և��;�G���Gsg{��M�J6ͥ��Q�grq5��(+�؀��ޟ&F�`�R䉇�k�)����I=�֖��Ǜ�3q�e�T��B�L�t�c�dnT�PD1A4��i* mLr4��\�*#t�>��N0<TF(�MZ\����������[�FݖK�潾j�MBe3 �č&��cV��x��!�Auqu4��4���\D��yh�y���a�6���#S�	���eq�ܡ:H~x�������b�ny��(t'7Hߌ�_��>O?_�A@�_U ���B��E��恅�JpP�&1�qp«��B����QPЊ{�S��������O[�mѵ8�`�=ٺc���#�{O~.	)������'?-�T)��ʞ̮�ќD�P|T�Z�7I\�[���$v���ВZ6�R���K�S%�����\ā|f�D�M��I9�$�n�1=(����Ɏk!�y{D������e������%����́��Ь�����E*��<����PRM�R20j�j2!�%��1i�9̌�jNI/��������i�j%��e���1�R��X�R*�k�� ��H�*a�	�e��̹�� Ж������4t�2�n�i���7R�~8��� {#~-(l��H�g ��`N&5I�sK�"�:��H���èpV��f�§X|1����~%a5��?m�y_�Mcp�m��z��1��q����m鋎��pk���ҝo�|8��sSW��Z�G�c�
�-@Y�joC�"4/�!�9�m7S�_���xC�A�J�n*UᎦu72����9Lq�jƦvH\K榰W�#�qQ<����F������1�d�b�����C��%	��S�������RL�ɤ	7	M&�"!��áдjSG@i��U�CB�S ~��y����G8�+��f�`�k�u��A�lB{dH���ȚkT��Q�`��Aqɦ�17J�dttč7kL�J6��48jv�i��7����ֻ,���!��0��?.:��F����w�&$��dM��i��8�&Yk\�Dj��S]��/d�
�y��Hܖ_� v��Vi�Ʃ���I����˦���r�ǩ��Y�OojCx��R{Զ	��!VG��]��4)�r���j�"P9��z�����gyI$6WX���eG-��0�-GT�n�8���d�Ӗ��F����f~r*���}M	�#\�	��f�		�#�����Ej�D�i��Jt�ݭ �%�F��SZ�j*�ӢNE���A�eۣO�:
��y� �p���b@�mA5�����b��L.�o��ʥ;�m���x�N<�X�EH=^��R�s��	ȭ�Vʤr �T�ּ�t�D�R6�%�4uО$�i�HOR�nޣM%��(hT�2�z��W�֑Y�!#��@�LL��>�����	���?�?T,-��P*R��������P���~O};���p�|��)�5N�pEb;U�̈�e#a�j*l,�����c�G͕EJ���@�o���6Zώ-2D`0t��ق8�P�y���R:���~6��[$F�(j�*l�F�� �̉� T�*{���M��϶��u1)����6~dm�\����|��t��ZT�D�]>�& �F������m� ��]��z�T�q�3˨j�\]-�]��Tb9���u1��	٦	�T�pꫳt�l�x�����R���&����Ne�>�<����R��4T�a�EQc .�:��T�e�+e��`�^�q~զa�P�)�J�č��Aa��0I1q���!�`��2��_hv~w�Z��ք��л@;ۧ�q!�jeT�%Wܴ����VS��ۣm���u�MAre��e�b$�Ҁ6����������luNW�7L>6��E��19i�i�ڂٗ�w�`LCe��ǕGcA�UV*�Q.���M��S��a<b��az�ȀP7**w̜vj�;5O܌�����j�8��(�-j�����ק�HOmy���׶�i�ɵ#S����4j��Dj"5)�e;jh0F���#HĖ�~�}N$sP >R7J�G�K#�4�h�^ZHmmKI���L�b~T�l��� ki�&�U$	@Il�b�l�b��pn��&/�ϒIū&��l�N�Z�}?yl=T
JM�wdkt��NLS����K&�J��^�0kڤ�"�2kdM�j������9M�@�_��e��]�l�NAsAB�x~�V!ҖLM�iO	-�O�����ӈ�h�2�R �O�i�����B��h���v�}NF��D�O��Jrk^ֈ�K7PIJ����I�A
n�-S�Rr���t*sy6
tŷ�y�2��v�i0��7$N-���ڍ�Fˁ��]�I�m�=�<�涱 ro�̒&7VCf�܄W_6�db�H�w++��"��Q����IAdD\�=H�)���2'��qꑫ?Dn�6�4�Ȁ^M�6ܲ�K_�F�f 4C�Cӛ	��!�����̼��J���bm����ea�)���~���/�}.�\Z(���8�nڪ�T�!#�9�4��#n֍�M�����i��`�)G_U>����ӒFGp2A�T*���~Y�z����Ȟ��uUN��DmO^Z�!�LyS���֒
p�w�?>�������dn	ж:�Y/�d��d�V:1l�D�M$n���J �C��Mʹ�m����bC-i�:5�j��}�?/PB}�F�OkL�K��i"�ؤM7+'�^n�,��G��ǀl�5W:��n�%��H��&��Ȍ�䀃=�d�28R��9�Mqi���E�a���;�)�i���ѩ���4�NP ��א5V%%�=�R�O;
S�R7i���NI��2�=�`K?mKH�������S�&��&�

����D�j�i���W�d���m����U�`���R�ャn�`�����0ml5AL�nl#NA��MAqRz�t��P~�KV�P����l6�?��Q0F�4�0t7[���MpV�n��h�R�h�+(P8��9�H�]T�&@Dqr����{s d��!A�6��.��Gd͠2�fO U9P0N[LvJR;���!�C*.�e+�T#����*��V�dt�ʃ�v�'2&�������y��`x����Hk����T���:|��(~l4�8P	��0�P�4k���[&�ak�dkLb�g>�j$*��=[�5��i����i���zT����e�5Zokbf�J�-��=���/���Rh�Rn}J���6 xtaEA��[}F��s{bUGr[sb\0��D����1��Њ��Z�%���s�J�3M@b���ZS�Ӗ�'��? �G8��r(L�tN0��9��S�L0��R�sud�8<6qH�R��U��֒�SD�3�0������Ę6�%�,I�	"c^KH���jȲܚ��#�bRz����914wn]y=ޤ!;�Au!��ޕ�v�j�kƫ�-jm%�M%$�d��mF�"�	 K	/������۷�7L��'��$��kS$u�(>!�ͤ��Ni	gg��OqM� Б!����by�`k�������0����eu�p�k5�^7cn�!,�e�(��<N���F۴�Dہ5kK1�{B�4�X8�ֽ=E<��Q��Q.�hTp�S �NvD�-�*�H��!M?�[~LvD�]1�P�4���ѵ�M�SS[���r Ok�̴��zZ�;�J��QҰ���:
颢[��A��$� F��7�վZ��D#T�14������|<|گ�ՙ,$�R�\B#Q�.�D@N15�KUB�� �V樨Ŀ4S�O[U���`�V},�6�5��]d�či	�WY>6
�n��N��x���b��㖫ئ�ll$Y6�-�v�iRL��OX��7�{�&��������h���{�9��6�&,��F����AОq�P�N#��� s~p4��@cU�O<��(@��s�=�T��I<�<���J�*&) �cYݭ0�]�O:�NCY��W����S����a�KR6�#�{U�S�Se�q�j�d�o21O�&��; Vn�Q�4���q� �#|���A޾yV w���3h�{0{8`*���B��%~oZ�ƒ5:@�mu��I�K�x��Cf�Q��e1�b��W&�I�ɕ�c��ǂ�D�0I�R�|�M�ܨSu�d���D��$N"S�����"'7zc��<����{HROY�#,��� :��I4�ޮi�$ǷB}���~��1;�N��i���ᅩ�9\ʆ���K�kZP�z�-�N>J�?J��hj�.j�.Nv��ܓؠ�T~�<n�TZ�7l�7&����$n�>~�Mژ��V�h�a��=�m�涁�bF���Ȫ�m����z�C��b�잢<�-;6�ڧ�FOg��N2�=@��@J1���{D������� <�b��0J  '?#��@�)o�b��˾�h{�9���q睟���>�\�2��6���R�a������Ȁ�mD݂2�����N��hD�GJn���(�m=dZ0�����ףZA�GE'�2�r�d��@$Y#L@m�����I�w�7I	n��9��5o��Ȥbo��RA�� ��r"Gl7L�#��Xt!�Ѥj�uڃ�0�D�FL��o�Z�)SB�Y���٪|�D:	��T s*�Z��41B�%T1� £�T	�s�	�5ȯ�`��s���d�ڵJei���zj��V� ����At��X�Q��'�D���[��bN+,	F�sq&�N'[�W�����A��pm׃��
5���i]�iC�"Z�ޛ��.:����崨��P�c���A�D��� �:���)�+�C�
W��A���-� 8+�M�X�jM"0>u>�X:�%6�*L8&�-ʰ�Y�����)���� +��-+�B��?�jӡI\�)��sKxb4#%pwy��o�j"��<ך�P��L�6�D�]�S�����V<�WCn��,bk��L�f�r6���ӹ���$(hR�<yR�3ȐJqU�^������i�Ǟ̮ qِ��j�h�w���ye)�;e$ZMu��EW�Ƽ��ZF]d�j���e%9����)�L��@ȁ:۫��d��6����G����!�DkX�$�!�i�oI��	m��r7l��I�C�V�nI��4�Ϯc����`�Cm1���=tu�ؚ�p���@��Ji �Q�N���[^��:��`�X�,��J4�נ`�#N����B�#g�瑁X��ڥ�& 3s��y"��L`�U͗6\����I���!�#fr���v����%H��E��$��Yj���Zwf��mR!0MV����9�����t�����roH(��#�5�0O+��F���U�]�~`x�<a�Mȑl�MR�䫑����%�r&��;����[��jokS�"�F���t���j���CJ`d0��TU���2�`	������ɲ��V�8�PF��r{�n�`�t��#5	�#G �h* 1��@��2y�Rs$n�c�b)LH���ktmb�X��
C�P�|&(S��>��*i��.�2� �i��K�ڎ@��n���
s�j�D~��$�GvT&]m$�[z�*[�{�G�Pn�)���z�Hvo��c��H��jP�X�S�I�����|6�n]��hi�"i�1mΠ�i�O��`���k��%����"j	KT'����l��[!�K���(9�A������1+��9�հ�mF�$	������T"}=9a�Q�4Z�[n��g�[F�GAs��B�0b3��2�(ƅ�Pb�#� ���|��0P� ��R��#��e5�J �K�#�{P ��1�T�9���
O} �rJ����Ge�*c��lH�q��r��e���Qka�tw��s��u�d�*�y�<|un�9?J\<���F�I�	�'1&�����MA���y1(���=4�nM�y�l�6�P�P�*:�Q"Z� �e��-M��Ć�퇩��6ڝ5c̧(=Z�i=�H'	�QE5S�۠��'� ��~2�`���ء8(cA�G��U"�].]���*z�W$�@�ꐪ�k��Phb�ʐ8�p f
2�e-c�"GG�.�@<&-��#��|���H�N��G�z"�)�������@�Z����0��"@KZ����kx����H�j@���Q>f�&���#qo����0�D�[u`��V��ʌ�!���x8��C����(�����G���y��5,�%6�P�<[�м�K�ʌ�nB1��-�F���KF��%>K����p��%�еjj%�Rx��5+�Z&7!r̆�p����,тҙ�7/��Ro�hD�kB�I��ֈ������_jr���w4
O�n�$�X��<I���-XJ#��5fq�m(!8�PI&��ޒT�l�.��IZ.A+CBA�S+�6\�7\�� R���&��� W��uȜ�����6o�\�<�\
Rst����=�-51��Lhy�[n��ګ�1��H�A��#t#T��e����đ�@�蜚 ��;���@i�.^7'X;��)�,�'Ɔ�图۠�'yr#���gu��Hu����S�T�m��@���H��ȵ8�_��J4���1�J4��y���o �Ф���ڠ�[ �ek�L��� �!_�^��,S��A�
���t��[o��4��g��nBav�*��N]3� hz��?{D	zV��#Tdv&^� t-~:�boe��6ρ@!�
8�.�>�#����qC��#�TV&|z��H�z�#O��9#��@=S��ә`����Qit�`��7hp�˪! X<����R���k�$O%&��ǝ�Έ�h��h�/́��O��o���9���3֖��F��ɵ-w�\D�$����8���׷@�M�P�y����e~�(��*y�E!��x��#�<�y�0�cU꜠H	@I�0�8 �cnϤ@�҅�Xl����cM��}��hi��T�b4Rp�4��y��DT�7sn�Op���c�֔&,��
č�ih#d��<~b$i��IƢ&�L�ܦ<|ה&;��2B72F��RsCU���s�S��>����Wd�'�T��ó�[�꓃Zos�S��7\�l�44ڣdOi]��L�1�H��Z �q�-33��Ǩ쪠]�b����NQρ>��"s={T��sPn�'NX�ÏiQ��9�_S
&֫T������u��>NG{8\1����!]a�j�.\������R;D��B)Ɔ������1�s����r�s'�kbGӯh�ty��lQ�ܺ%G&4Ӛ��s-4E'�[F�R���N$vrY?)��/�7�E��c����*<����qBܠ!]��i�" �:�K~l
)�$k�f�*6��cgGtŶ�Ðc�B7b�� �TZ�kZ���Sʚ�R�����]��eA�0����Mʊ�C,�h\���E�˙�32^�s�B+E��U\��� ���FU=�-�4ӑ��ҹ�� �2d̹��d�e"q4��b5_\�m�M16�ɯ��ݔ�A�b��.[;�[�i�H�`NS �ķ�ZO&�B*�*���I0���6��Z6+t���[�u|9Q�ρqZ� P�^�x��:���h	��p�(��&�Q�%kh����B���uM(Z
Gh|����1������/%57���^p�h4#w���o�:�����Zo�~
�x��1q�y��s���n��f�U�A�xJjD3<1�ă�8X8[B��v�l#�Ț��vQ$[�~��e�e�l7�$ƴ���;��M�9iE*�*��h����Ҝ<� bW�O���	�[^z�q�a������B �;ulCu�x�t��{p	���@+��M>�-
r�
���Z�8�G-Y��^@�@�
����I�i�#rc|�ډR�o��f'C�"BH��/$����&')K'OYh!�A�Nԣ��F�A�Ȁ#d�����kޢ����z$�ލ�)��$h���5\��N���	,�
�6�J��1��0�����w�u|L7FA��<���7�D�D�i��\@�v�PK=P�Dki�[��Ġ^<q�������m$�>ȑҏ;z�\��`�@���[F�V�75�ؤj۲���@(&K�b�{��k��`H�R�2Z�n�������ґ'
w�6M�i��D��"a#a���ӧg����غ΀6�5�q�W:�	V����6�s�ZQB��2�O���c̀�`�ndh7Z#2ӏT����&�7-�A���4�(&�����@��"�f��$�kV&�:��DL�z�4���=~`�[{lSۨ(&"Nl��$�{"�:)�tSU$�kD�ǜ�����-Y&	����9:��%�'ԧF�"Y"`��ڕ>���k��Ch�H��+D��ceE1��i{^n����l�z��shI6��KebFɉDm#_��k'��m��j� OJ&쉪���V�+U���>�����������l�49�S�Z����umsu�q8���t���.y����s�ǟ���1��� ���f��A���B�&���Q�ȡ�g�����" ��8��r:&�p�wb�ϥˆ=U���(F���W\�/���{J�:��tE�L�.�V��(iP~O{0(S��Gs`�4;�]l�*\~�)�$�i���H�*���F#�{ �p��$�7�H��%��G��;)�T�������{@������
�e�$N�E���m"�["M�#w7����|�2n�s8�F��4܏9`�>_�#Z����ڏSF��*UJ� {?i��S�&n��>i����E��~O0vj��<�

�*2��P�#���92)P��OPh��TЂ䨚�\]�P���i�l��-�>�J������	C@d�j<�rX�7N$R[$i�yYN�W^(�S��RZ<�u�Z�j�F5�$�&Ԗ�|<�M|d6��|�#�_�\!���8�^өZ���"u����<u"?�q�*�1�����(��x����� V���3F�ja587�,�/��)1�x� W�x�K���V7���׋Aq�Q�H��J�:��\��d6Ҭ|�5᎑Z+�BM��!i��L5���V�ku7� ���pH��5�&d"[ 6C#D��#��E���t�ܟ5�Չ]�nڛ�U�j�<Q�2���e�]�h�UesC@��s!��eS�f� W'��2�q'�\�N{�r��y9��l��� a��@�����j�FH�e5j��8&��<|�3�i����sL�!M��kI%A�Z�h���n��&���j����g�&��I�$M-ki�����e~�d�D:�JF�J&���(sI	�"Oi��"�kZ��� Pk]���	n��C�O�v�e�ʑ�V�c���|)^�n��B �"�����r��F턉ݪ�&�y64ċ)$�PR�4�L��)$�����0P��f���rhn��G�&���r���׻F
]�ٶW(
��t
���n�iț"�s�ҥ��3慳Ә)ƙ��т�(�̨#�l#ݏQ�%Eȝ�&�"��^�ց����ӌ�(Nh"NL5	�@	��3c��T�'1��$�r1�"�*��Y��/O���2�ckAT���H�u"e�y��pE"	�����w����\�}#vs#vD�� ��]�F��.JC���c-S����DiR����M�`)���]hW������FJDd�'{��Fn�vj��i�vn���Q�#$gȎ6����¡��4G�C 7Q9i�,��,\܊�7j��F�Ư'Y8��}I6�}vOt(�P(2�u�ڕ�G� Ԑ٤�����O�"I'6��KKN����~@��}y#�[	I
��;[ ��h��O��?[\��	���r{���"lPJn�8�n�~NAp	w��L��e�D���~l
.�e� � 9?"Ў����ᖊ+C���B��V2�@b'��YvZ6�v�Q�IF4P�2��*EAu�8 ��Ԑ��10�1ٰ�)���Q�E(�?%@��*h8x�:S��s����|1k�|�l:�ZfQ5^�N�!Қ��~D�~hO�V�D)��TRV7'���n~^�8�`58�S��P'6��bp�e��RB��4T�'D5=�~�M6��f;���z4���mٲ�o�ef�.5z�Z�&���I	,^�Z���;U� ���&`�`��F��v~�<�T��A��.dQ�"D��p���4=����0AqV�R�h��Ty����eR��	@
2��)A8�ۚ�Q˴em�%�a�	���}t *D��6�� Nj{jSj�ɇ梱XD�6(�K[e�wG-_�O"Y[���%���j��kt�$!%�]�ו�F��zY5��@�'A4��SX�I�iMf�5���t��If�D��Ȩ��* kOȖF�BѶ��:�0$:#Z�ț|�n�}n��(?'�l�Vڮu�G#�Baz~:tN7I;&/�JCq�QB���:>�8��BE1ב0�H��$,�������ڝ��ryh��p0��SRcz�<P�e�	��nO!�kjOF�Nɍy���j�-�Be��4��UZT)Y2���]T��CN4s�|�~i�?4Ӏ6�Gc�<2+���hH��ֆk@��C�	"��хh���2*�_�4����y��Hl5.t��	�!�)��hoK�Q��e��@�S_ǚu9�a`S?x�M�J6�����ٸ)��{Z$�&��JD���BV���0K��U�H�(��h	7�j;H(�����)�274K!2%(��o��))#��2(jAX���2���4@�$|�׏S�#��w)wCf�z�P�r��I�ֽI��rʠ^3{h�o���	G_[��hb*>�OF���E\��ڪMXd-u��ӏOg��B���9%J�d�������^E5"Q���-=u��u�vUl&��Z)�N|�)��J���\yh{H�Wǅ$��.����T�k_�F��[_kܮ��Z4S���d����6����m����M-�v{z��� �h�NՌ��#�P۬{oO�	���h����(&��M�I���cr�G;����Ewb�9��}O�Fd��:~כ��\�	�J��s02�nd�l����oO�7�7"Y`�$(�n �P\�T�w��H����A8H���z��CW	��;6ME�F�zh����yд�T��s��t'96���ԩ����D��j�?N@�͂nl#[DF��MAQjr&���1�~�M����rND��r@�mqBy�6ɓɔ�G�q�O� �Щ�1=)u��S�iW\�R��~=]�ZҪ8��D�y8���n�~�O.�`��bx�#��QD01��bz{em�wぞ�#�hJ����V��K]� 76���aH�݅4
<�(�@�֊��yQ�t�<�����T�x����~�:"0}�E(,Q��8�w2�ϬЃ��	�o�W"�I��T��vY	�N��h>�$��LT�r����4.�`�v#n����j��ݥ�\��g�eo!�w�5HV;��	�G��ra�.L0X�S�����rDM��:'bCr���A�<$N1)��' 4j'��Y�6\�>��(]hc!T�S�CG��	lawփ����U���(�1Q�Ȍ��掠�e��衊� sLLL�>T&�r��^j.D<�
n�T�)��m�>q�&\M$�$ޑ5�"���MHM-z��ڮ�#�Tl�Z$b0,���ŗ�zOIJ�I"q"���#:�N�Jrh뼲P<mIG�CT�5 ۠��,�E�c�4Bt7�'�.�Y��H�W/��yhd��5I�����$j6���ӳ��vp��h�zD�q-	��Ěvp������۵䴋jKo�%�	�|B�6���Y֥e3�L�1�K�Ģ|��Ӣ���H�΍���rk�m���Ħsw����e`Hi'�j�;/Ĝ�g��tuԶ%T��T6�v~@1�c���K�@cD�����܌�C%�`||:Z�T٣�rx����׻�T���DSw��#czDNoA=L�D��y5Z�$Di͂���%-^�����j$p(�M�~Ӑ9^���Ԩ$ֹ�^G��fHI)0y��NRpZii�����U��8��}k���>l�0>D�P�V���\�2��2Ŵ/����\ ��8�n��B7L�^;*~b����?�KϕH��o� �)�"q�4�'������D�e�~ا�@�����;��$a��4D	������S��Qg&���ot�A�ݩe�xjl���b����kBsB;LbT�9%\�pMl#e��f	��-�z`��.�(51�Z>�~���i e �5$�WR9�@��zR�"U��0�Z��fъ&�1��R No�����fh�5Z\*`�Mї�-�(�b`:�7_�N;]����U�_T��2��L��);ߝm��DL�:i�@kX��ܘ6]ͭLDHp�4�q�wԓ�S^Z��F˼���%��v�O"s})��&��-Z���5(�f�L#48�����`�Z�6�7N��穱HH"w�D�N����y��jWa�R��ӔM3v����FP�5T��9^�[ -0֘j`)�S���`��ǹ��ӕ'�����	��>i�i��������uOuOs�75��E(#�N.���1���F�U�.�n��E MFO;[j�6K[���bVq��"��~.�(!A
�S+��h�0��1�w�9�4#�4
<p�E� e.��
�H.T�,3\	P��Njp����ݶ-�ʛ���!�	�� 	�dm��Բ���h�I���3���F�=Zc �kk��S|�0t	�?{������'&( ?sH���*P4��
��h�M$DF�w��ͪ��jY,\����N͂"���Bi~�����h�I�sy	�P '5����ז�ͥS���r���0c�
;E�B��W ƃˎJ\1�!��?Te���v��U�䨐8��	�R��������0�H�Ib�G�yɦ\��ۤ]�E��Q�Ct���dt�4���DM���퓸�����-��ґZV�����F3x�|��Siu>�Z�q&�$���"�V��SRQ<���\u��J�?m��X��%V4a�Tf��W�䋬q|50�(�$�mI&CjO�(&CjJ��оy���SS��F�cqHZ���,���x?��*0��n�CĚێM
��KR��F'kȜ�V&�bĲܦ�jV����Nū4�ܦ�o�r�O,�R��*ɭh4�KW��5j��"�rkI�CU1i���6jkM�ٲ�M*L7�=�j�����Ю�J�rA+�U��C�t�HhJ�fyu�'�f�uPdr�
�HǗ�R�27��g3t�6�9������ĒOm]���i�DiI� |\�=�m��6�*4��/���7P\�vMw����jWzz�4�呸�A�t��6_�F䪔��4s�2G���+T����bDdFqHFn"56ZՓ��!��$�  Pn~�yyϞ���5`N �-��]��E���������y�D���[�������U��n��F���F����4�橓��I������[X���?$�ݞC�ǐ.���og������D�N!�bh�ɯ��0}#5=^D����*b{E���g?�S��ZѴ����ջ*}���1�U�TVs~A��у���pũ��(7AJ�¦�t�er��yeb@S_�*90D�״�7��4*G���w?��Q�i�v0}���9���j��W�����'%2�3T���MS�5��֣J�ӟg�ʛ*kl T\L�D@MvS�ܚ�t�L�HP"z�5��D��.��֙��l�^�(��D~��T��Pa )@�呺sj:�jF�TD��k�,y�y#�����ɦ6hp��P0��J;,ۋx�!=J	�k+^�;�*0h8Pq��A���sH�p�P��q1���';&-�H�-�U;>܁[��7\���j����Lv�_i��>NTn�2���Ͱ��~�S���O�Qܞ��-�4���~PT��;��H�iZ�Z(
A��#�����b{�cN��L�U�]9�a�L���(l�.����@`�4/n`��
J�TJ�na���շ�N@�+o���*��44[C*��"h<�Q��Bg�R��'����ǉjp�;�+`�l�٢�3i��V��(��V�)��$-�����#��ȡ�ޒ&$� '@![h��q8R�kd2{� 7}26����V���#elMtI=N�'#���ؘ���Nob%�E�Z��JbY ��YW)��2u�( ��� ܔ[�&*$-�-��T�P~�(D�*q���eR�*h�U�eRV%.����-v��E��bTT��0� �?" ���(cJ��Au�9�B��o�l��J�l�I�B����]c��n�_���"@�Q�C�~ެ����2�D.�n!v�7)0� Jm*W�|H53�hNR���_�[���':�CT��ڳ;��)p���8t�c��J���'+�a��n0sF�%��R_<�Ea��-I�!�ͺ1���ԔԒ+A���M#q��v�����1-�u)�a�x9|��`�Ni��f9yԮ�kr�I�����ۣN�����6MH��Ve���^$��V��kmZ׳a]�p��J��qi����-R��[�S���t?_�+�UNe�4%�4.تxQ��W�S��?��.���Ј��#��g�NO��V��`���S��G��S�c#[)���j���� P���"#N� eH&@���k^���@�K!��iI���P�W�$�j��t$��@�`�n��Nw�=���-s@�8~�֛�|`ީ݈�6�
� ����'O�M�1ʈ���F-��	�*�ٹ5H��ӗ$V�Wҳ���SWc�6�hF������$$
!-P��~kmHۓ��r�ȤP��iH�pM,T�f��fs�J㢅�T�6Z*����xQC��ĈM� PI$[���N[)n{��Gb����7l������6���F�rhx�Br��ei��
��rV�d� ���o�
�[���6��Nl�����r��ӏ��g�������{EQy㚨d�w��BkpY��T�0mI�&�@"B76��i�Z��>���ѭ���l|�]H�HkY���Ҧ�eɄFI�,�m��-��m�K������N&��(6��o�REv�4�+�eq⒝qR9�^P�$�7h7;��ě�y�a4|��[vz����.���!�TI���ᖚ	KN
t'9��J	��˜�l��`�턮Iȓ�\����l6R�['��'�.j�l�4?
���n���>h6��O#�:}ݪ(ښ#y� 8^����-N}l��m�� ʆ9?4��� q��ǅT0�#Q�'?%}J�v"�@%MmҮ.��GJ`FZ�M8کӖ�ӔTG��euu����v�QG����QhR�9CeB�45Z�TQ�c�N�z�y��X��2����̹%\��`�=,V�9bP:MS��k�h�
���1N��y��5���#���*��'��<���`�rz�#P<�?-��v��{����Vվl/��ɧP|������berͪ��ޚ�������,��йMa�1l����+���`4���~���K��.Jq��uʎ �H1&Q!�CE��<�g'����*�^{8��e=�r`|nk5���ד����r�;+����ڬ%�h�H��'<rb�馔���"MW6�L�&��9���$B�G5���JC_OC�
��c��8��Exڦ~i�Aw
1G�[@A�-�1xCQ��#hZ��t��\uZ��"�+p#�"�$V��󯎧��-;�D0���mDO�ո�]c���84��#�G8����(&ۃ�Gg�RH��R�鬄O8�|�4��D�	�д17$6���_���m�5�ۺ���L�OD�X�����L��޷Ċc[L�Kl��"���F�����hf���O���#�<�qr��J��?���Q{B$4*qQ���� q�����ҽ�@c@&��5�<� (i�	��.i"KU��rP�kt���B5�xu��5;��-��ev��q6T�W%1��DR �+]�D��#��]N(�D���D�s0+/��N�S�B5m�~~]$�F��Q���S��!A������W�~<֩�7S�8��1�ݲ~�$���-���d�6	�d�bͺ]ٵ�?\�[/�	�#ճ�
B(�ePL�څ�@ȥ9C�5$���\$��f��L�VJՀ��}U�o�oȞ��h��A�g�T˴�NW=[�+uٰ��i����B&��<���T�n�(.T
g~�LG���if���6��dɻ�V��D�n���>1:���֜����|D�+���S��u��rDr�䞃��ޝj�J@�"~�Oy4��n�b����D����~[v=h�j�x��Ę�D�rsGi�Y5�m6�c���G2҇�҇�q7��E������?8@����N}M(H�&D�9ݳ'�"(@�&�Fۨ�w���|DVS�Jk"k|:ww��O�9�?GJ�8�S�RDĐ�LlQ�U�bb#%��ܕ(W��!%#T�Imش�	����%��1E�[��Zg ���m��T������v}��Zm��dN�'U�M�����t�f��J�R��J4�}������j�5C 	�i�g�����	��rǏ=�J�f�f���Dd�r*-(�.ɝ�2��<(�V���a���`&�F�G�֨�
�*\]s@���Ҋ9B)�3���)l�\��fȠ@*��sUG?vl�ʣ3�&�ԑ���H�����g��:5=�$Z	�n��i�A&0�5ɢ�^�	����TG���@0��!�����23������kt�ħ>��[�DOSq2q�.�o����i�N58A$�r�T�{A��ԑ؜$ioQ��1�ܺ����X��(~J���0��ԭH���*�h���r��R�GTpʣ�O<��Hl�h�[C'�hGJĨ�����(2|�l���T�!P"hԩj�a�� I�-�I<��Okەᵹ^�� 2r���nv�"֬���^7���+Aq"��nĮ�jn��RH-���I�r4?�`�9�VC�Z��V��e<Hm�|���Z�r�p�@�R�(��|�ngY�%"�P�h)��͉��p��U#j�6��u2�j�1�N�~�$ޛp��_�Lg����������,����\HBo��/!�4�hg�p^�Hj1�jC6��B����m�@�u��2�n�*?�9>���u0�	f@K60w�(�B���*�"J�]��S���Xy�-�˗�p eC"2yQ���@�4.T0��B�@cC򃱀�@"�[�e&��v%�M-6��[v.��AAbH	�Z`bI[#���rD��u��ÃT�i)`�D�����i�o+���5_�O}S�=[r�٨zP
P���ɦ���`�aqk�1���a��`�Aw1T-֫d���㘤Ko��tq&��hMf�խ{�LT:��q�ڣ�I�F�e���w6	��Wٻꢧ:�{�%���"s�fw{H��)�Z5m)�z<�\:����љ�v2y��r�r�z*�l�����i�K��e�d��%3�Z̷C@"hsT]�1���9Q���ƙ�Š�ʭ��FѵD
���W%���^�+�kQ��7�@*�[�������M�)d�vj�	nfã����S�M8ڃ|T�X�Qʟ��Uv�" ��(.D�A)�����l�?'�i����94P2�kǜ�!���;
l��7D���mi��@T�l��[��	��洴����I�<��*'�o��J����"0K{�x�~Y��ۗ�:���a(�`H��ڏ�W����|F�$�:��������̑�1@g�0	�$��I#��� &�9/ӎF*�2��it����5�� M��=_Qԉ���2G4s�.EA��Sۦ]�k`��f'*7NT�}�[�k��g�����D�
�6����e��b��ĥ5%P�l Z&�����98����Zbm6�!���@��D�Z4,h]hED�R��.����� D�e��� �����g��̀n������92�]Ͳ�����a�C(�%Dq��`@���q�)l١sl95H��'?(�=J�2��V�d��״W�P"r2e��d�AmbH�thP�]�b�ث�Z�L��Ib�s-n�@ȗ4ߌ��.���+�&�ԡ�M�3���Sƫ6ܚ�oED�kMH$SM7���"�e8�Xj�H��w��d
bb�JOG"?.~�k�#k$�������O����A�rR�~�*���2qQ���.p�v!b!��j�� �TV�p�$yu��ϝ�H�E���E���M!��I8D"Ttmm3s�a���v_�ԥ%b���n%�$����R��q�) p� �ԩ6��F�C �y��#�q1�zL�"�)�Hm��Fƅ��鷋ƦjJם�����_7�\�����D�:��"L_�^v��V��6�
�o �a�K�F�h�^�����z�N�A��mN�Ba��ln[���xu6�i,.���i=DWX��
đ�f�%�Z�cHm)$	�ǈI"J5������'����A�ŠB���	�	MU!�ԦW������m�d�~����C??=�J�/B�K�*�NJ�S���g��s(��.8yʨ�hcB:U�G<]��Q��U@�rr��tt����A�Su8u�� M�����G"O{I
5	"Y	����we1�=�'.6�����GH���ZM?/���9đ8�nG����0
��ӓDH�ɔ�#4��"{2���T�옷~< ��T޽VEsK�Dt'�U��#��9Ca�z�W_�#.c��mU�E+M���#�ݒ�a�2n�n�T6�.�#�FZg7�G�3H jj��6 �9�K� �ѻ<~
��*�ĮG���i��z	���ٚ������������>��q��B5n�.d��Q���| ����#hy5\���u���7}<F��Yw�$C��{�r�5w��@%��V�y�SV�D�Jd��Q�䤊r7�z=�b��a����ep%M�D�wyQ�H���T�t���g����Lrw�9-�(�o���j:]s��8�&`ܯ�6����D���x�h�cAA4�֧&��VF	�!�h54�֣dnl"vJ<�n�����u4F(��ဧ�G% 5����޶$554��C��������G�v�eH��n�&��ҁ��H�Ҫi�Gi�rA���[D�l��=�߭�S����it��u�Îf�ώV�+uH�BV���_���>��9*}sD���UȻ�L��+��1�t�����PT����ǕY�Esi��s�eS9�UOGh}J�SBq�xg'�%Dp��c��E��~J���D$F�|�T0�#��?�1���n`��hQ4.��D��"BЕ!=�� >r"PP�K��N3}Tq��)���ؐ�)CM)�⦝���J�0��K����0 j���D����jy��:ںk򅱳�s�dM�MՐځ�HL�YHH��1Jr3�����j���(�|�k]�S���ڌI#J���Hl�V-6����!��y�R'5Z 
h )<�����A�R�*�PapOh%=\��$G��.�)�G��8r��Z-��TG�\�<(�C�ɔP	E����	��E��mU�H4�����*I���\m���R *.�#OF���u�Z�:�~��<���J�<�H�T޶Hͩ�m�t��{i���$oRhHD`:m}Pz�}#.�:���Ū��{2�&�cV��~T�vPGD)���u(�*i��ȹt��s�deBI�g���0����bn`�i��O�&���p4��2ש���:9�����F�fѴ�ԍ�VL Mn� �ٴ�evq���׷)u�ҥ�T�INé"��W{|KR���Km���+� �r!�JzyR�q���'�]��%hD�����FU.�S��.a�7S�9�~>N?X�����v�~ L��a��}�����b+�����٢�*sT&�1�'z�mi!�K�u Bn���u3j�)$�;�g��I�����T�-J�~mQ�MY$�́BG���Bˠ� �Ct�l�8��e�� F_D��ד�#d���@��F��Ђ�z�GJn�r.e��~D~�#j��"�Ր�&����kdP�AQQH�e~`bG>��~0����`��!5)�� �OKGd�рEs=K�A��m�D���e,�=�bZe�^����U�ͣc�r\�_�=��K�7�����<Zr[��ۚh��������m����M�����!-��K��K�1��ˠ�� �`��@��l��(�������e���R��B'4H�e�mZ>�}j�ER�
hL�P��@�1�d�$|�kJ��&���b�K���ɲ1��~Y6d�.I�!� ��[DSj�!�fE����Ar�E6��'&�hs\<�0/*1bn�ڍ�I5_���h�e�"F�mm��l�j�v$}{F�svD��r�#~[oL&$kڝ�-3O��
Lp7O����T�C�m����X�||�&)r�}��K[�ک�A����d� �r�����¢D��[޷&�@YGL<�)��Ěm	nkj�fL��s<]�R$vWk�쥰b��õ��� ����.<�͚�0�4QУ�G�'����r2��O>��B�1�P��[E��.��2�Ʃ!h&��@c*�bTH]]{rvl�Z��bTr�A�q�Q*а�s38�G$kD�7Q�J�V�ʝ�o"�M�˚`�B������P0���`E���Qjp�Bq��t���TT�~�*I<�������=�#P*Y�,F��9\�66��E'Ӻ�$��m*'&���4��=2j�L���QSa0ڧ.$E*n�����@ndbb����ᴓ����e�Z�<����&OP� y�R��3hUA4.h<�K�A��Q2�]����S4 �y�����h���26`��=_��SjJ�}-��b!�'x��zޜp)�R�D�U�' �#tmN�)��&��7 �zR,�'�s���$�N��Mj�)+�kU��|�'+��eJ:t+����Jr`�<u�$oB�m�8uHKR����8�uN5 Y���b5�V$p�I����Ii&�Dڕ��'���  �T�1@4|�Tv����V+�*W����-F�����G%����[���7Z�����-L�,���F�ȉ�жգ�A���$/�`���Ÿ�6��Loe#�DѨ�k5��k��!��1q�������K�.m��9͡�R$*\p�R+C8�S�įc9�����3�Su��_�����HajcB{�B{��똪�X�BR��}l���� X�k�����v����DóZzo�9$�$�G l"$N@�y$Z�HZ�VAbնR����H����~#l�7O��\�)lM0�N$�H`�|��w�������'���F�`e����đ�I����!�⦜R�1�Z�'�5\�5V�-[�-[oD�6V�#��������9��YS�]�Fb�LRyJ��{���[{G�L�
�����"7&��k���j��ǵK�g�U�j�*�����4W4W�%���F���ܕ$i�i�.G���	��e�/��$�;B��6�*"[~l7{��\���M��8:��$�T�/��m��g©�Cf >ݏP �z0���@"�`��᪓�pt�4JH�L\��T��ٽ@��ɺ]d��5[t���i���)M��k�z�7$��W�J���sѰM2�T.�r5�oH��ۨ��j�S6��-NoG�k�������$��$�?Y� �?L�	�Ԇ � e���'6ʐ���"Lw���eGS� 5�i&�۽@�N|�X�=W�Q��!��@$i{��"S��V&��Oi��풧��7���ces?
~�Hi0$NDz��8�eD���3�9�� xa���V�v�-
���r%�Y��ZWW 8���~��:�sF�Q9s*l����j�i�oϥ̿4(5V�>��vGG[]�RW�����;��qu��� On����Q1ʌ�#�2\�#̴U
]U�X�yl����]�3(�kh&#�-nޏ6IOܯ� ���2��0�aHhT�'gԫn@�����<u}d���mG�� � �N��-mW�g@4�	�"5<�	&-�^��Q��K!��9��Hj�X$L@�8��A$<~�p'�ǜǑ�`Tr���dE�P3��R�n��'�O.�h�UB�'�9�Q yc4PED���l�됮�k��W*cA�G��Tqu*9?1��pt��$6	H$0t���� t3�PU$N:Oͦ��g�%�ţnȉ��Mޭk`��6�Ձ%sS_�֦%���Z)��58I�:YXR d�c^kZ��r�d"_N��]�ښee�9I������:����Kq>
����vI�Jm�X��!6��bz��)4� j��W�KRp��o�ғe���r	T9 PF�{7i����SDk�����mMQ�� �&���E~iZ��9M �,�W��~jY���à� `�;�P(8	�T+h���`É��2��h����	ѵ��454���_V�eR����BЩR8���˽�"2z� yR� qr#*�<xr����9��X|�xL���2��n�{(j�*j�4���Q��#{Ea��	Ǐ�kg-����O����4�<����Њ�$l,��6' ӎ��5��4sU���]�)��gE�0���<`�(M��<T�:�.�vP$0*I'6W�EڮE��� :
�y@4�-shj�"P8:�pJ�Ӻ��U:�^���}n��%��ˣO�(TTڠ�7i˦�{��eH|\I9��*J~
q�Z�n��m���0���ڭk�����OT�7c�2�K=T��U�GD��?"���(Z����`��b@�5C]�-�*}h��m��}m+��t�e��4�̎�[��%��%�X��NE?{~N?z�9���2s3\&������@2�Oȭ�H>�=���A�j$��
7[>(|�����w���	9#�<�GLT�H��Ml�6<�4���E���mb�DDe�M#Y#	bN�������$DƵ��e�:-�k���C��rӊu#J5�Nw�kJ���� i�����{zP��j�&鉢�%��i��W{eN|��eP�� 7#���f�L��1�H|�mGM�E��  � D�4�r,��G�J�F�2%!���&6�~n)�Z�IA�֎�@eM�P�7�ͅ˃fa��F&<�<\��4�l�L N[j���P%ǆK�cB=z�t@�(��}3E��V���&Y��h]T�t�2&�"&�p���4�q����QhK�J]������cF.�\�ꋻ?s<�)�G��������q�A�q�UZ�V�`�`��n�����(&�\��H�����#�k�Ț|E�*9�s��x��`�'�7Lb� �MW4h�����)�[Q+���F��-$:���xL"4�Ȏ�� 4�y�L: w���H�l�6�<�jѩ�#Ry��y�n	��}_��7PT|�F�?l�Nsl#H�W��2%N`��H���̞A����
r} ��<�*8�4*���H.]A
�\���b�v��TG�\������Ҡ��{�=����������ч-6��aL0LkLF�Ѫ{��G?>z���K(�����jhu���8حS�T�$�p1�fՂ���kT�f���l��Y5f�
ΧA��$�4ܚ���ݾ!�����H�k5
�u~V>pQ�@�#^O(I���k��n�)��\Cb��l[LRK����K"j@�u�N�đ5 �)/�楃��j|$MM
��Ǒ�`��А:���*R��FǑMxj;�R�ЦہM&����.]�<1=��T	u�Jҧ�y�h�vR�m26��4=M����h��mLI%rO��6��(iO�yb$�h\ƅ�h]D�IZh@��.hGJp;C�JfKS�]��`ȫ`�Pr���^�o���.v �a�̜E �족K���A�*ޑ�ʜE71��=�^�%(ԐD�(7u9y��Hal%�
~ ?D�~"L.Z�rw�,����HjР��3U<�t�e���{\P���$l�r&��>������X�(8	4��}���E�l=��V�^�[��#��<ԉ�e�|ZNX�y&H�^����u�7�F_r2�n��-���/̦ ����%��4��H�ӅC"��7�
7{~F��J�=�l�T�')��s+c*��"��j�n���ih�MW���G�/����#O�����ET܎S�̶@ 	�ў�0�x�#����I�"��B�Q�ڥݞ�G	E;�f�A^�n���:�dM��֘&�I̚�T�lȋ�0\��hT^3~�J`f�%���O�n�
-J�%�,��Hڿ���ղ��{~}{h0\�)'���)ʔ�o�kVD2~���F�m#5?�������NoJ�'Zk�5H#�h����L=i�8@�(7<�4�D�l4/�ҍ�Zk���G#�5d��>2�e��<��:	���+��<�����@��9�q�^�\����'�eOf�#�������J�T��=��<�4����
�K�h�qvZ*�.h~T��&�+��TЂ&W �H�A(!T�V�* #��44ߋ���&�iX�:��
{��Eh.�"�PT�e+�<�*��(�"��{~�"hG2�a��]U�1l�b<]��=<x�aS����k�"��3��~ܘ�=[��׵!@������mT�4�t�1�����P}L�=���,W����M4�RK��i~`"k��l�:��"M�R�$U;�ֽ����&�Ѝi�z�SN���!\��)�j��4��p�#�rvN-7~� |� n~q�� * RW TW��&��#���i�i_�^�uU.\�ЉR���8��1V�]���%D����Q\�ʩ�UZ:���b��ntH��',SO�� 2a])�#C`��@�m�$3�IaT�H�&�b�S����m��dhoA5fCm\I���SQ:	���=ZjnG+r�ԑYՋ"�H�k�jsR��@Yl	\����Ҁ�xڦX��D��jZ�)9�5�e��t�&�!:	�ՐIHiZ�	΅d�5�r0:5泠5ֲ!/+1��"bm�rʘr�HSl�]&��۷���Ė����bթ���m�xIHRx�m�NLp�M����&��&$�I���b��2��16�;�ȒC��0��5�i�5�#�C��{U ���-��@���`Kf�*�EeʚDqu����heP$t��&�!��ލ57�c��a�'��Ll�� ��:F����P.�
yr�I_�.j��fSCn���|���7&$�A�8D������)
�7���ˠ��~5t>�RQ�	��	���R��$7J�N}0?p�(n��6L��fn�m� ���I��fRNo���U�g/��2�i���ѳ'y��Mt��d��.�
�f�TW1"oH��� �&�jG"~8ޛʑ�Ǘ;�����_�\u�#����ʜu�D�@���w�둔����	rS������t��@ʜ�q�x�V��)�r���T<���<��
������(�m��LP/N/}= ��1�M��F�hr3~������h�#���5��\��c||:Sj��m����������&~�D�J�i�5	#W�#��1�j�_�@�|�n�#?K*OEn�Pw�E6O=�O����c|TY"}oS���:���ӻT��do��645�5��4�f�i(�
[;��ZA�ɷ5 p&4ͣ���BQ$��ʑ�o� i�jC��`-�*Z�P*� }A$ӽ\��S�e�{�k����Mr�f�.T����&
i�#��@6
�#�_���}�n�F�0p���Dj��%�/�Kh�>�P2�R�W��(崙�L�D�	)��L9@�)uS��?�1*UȐ���ʥ�UJ�v��)�$�NP}G�J�'�T�F����M�N2���m�=��h� �����g'���H..��Uu90l��1�Su���*Oz��h�S�	�#�[�6�ym� J�?��ȟf��'�L�� �0l8Ӊ�FP�1L ٸ���jĖ�n@6]Mӣ���;'��% d�A�6� ]4�S��PBMS��!5��Un�'7�����m�i�'O�T܈Xb籇�%r�z�?&Uoh�`�� ��E< ���Z�0A��g�U"�A��1$.D�Q�ǒ�J�r�X�he���O!<�#��J��ʭ��.�pc*�?U!h\�F:�y)�G��`n�G�f�u�hrL:ZS�G@j����sc�zSq�M�j�m
B���I��M�&�����o��n�+$��f�,��""�=֠Zޣ�����Kվ4$�������d��Nl	��e2 5~כ@ԛZMH>�%a��V���ؘ<V_�V	���$MH7�t�9"%�H`m��0�kzSi�[��x�4�6�����;�J9Yf9'���3�Z'��u�0?%�ևBcHBR�M���)�*CH�bw}L'�*W
�K5��M!)�b6/�F�E�4��I�=T�G�!CE@����Ȏ%�D��MY���.2���Ӂ�����69>�s{ ��}j�Q9��\��}{}({7j�"�T�T`y�U����t��.���ֻ����ɇ�'Ah5�l�K�E&����a�Jَ��7�m��^1� �^�&6�b�[ ��˵S��T�n�֫LHM@����cu�1���8���8Sa$6<Mk^�-�i�n�����˵S��'�6@6V#i�!�D�*���#^C�Zo���VH�ʘ#����M�ѡ�mz�"����fn�<�2Q�������Q�W`�_OR�j��������q�xR�fT��Tگ�$�&���/m�"�E���I��E[�Wb�����j],�k�cw'���)��${��p��kt�d� �l��w�"P�~p4�BT�ԯj�>��S7�������8�|گ˵�l;�M�d�7�-lA*A��l�����k|TM_�F�\���w&-�O�Sπ�����;,����%��Cb1:��l�bSRb#��$�b<*H)�Nz�M�G�9��Ѝ}~_��-Ѡ�o�h"��ִ�˽>`^|���۲I19�s5�S�dH랫nm��0��%ͅ�Q�օ��'��tH�Nwd�OnH�����������'� �Ȁ6'�;4ȓ�5@.}B�<���(2`�+m
�ND	=ͦ�Ï˟�%�\��B"�T)t�]��	�H%\��r%ʑ1&"Ef�U@����
��e�VN"�Tƅ��Q4Q%�{/K�N9� ��8����a�CU�Z~~P`�j�r}��]��Ј˘e6�L��ʃ��c ��܄��i"&�j$p�>�8q��ޑ�I
o��o���S�v���i�y��*T��-1) �*Nt����������L?��a&���ڌR"[�?�=Ӓ��ѭ���Y#mT�e3��.Yvy��
$�!���ڻڧwC�����ٻ�x�~Hn�w����dB���۳*��s�Y��h�b��Ӝߜ�ZW!\�( �H�\�����V�H�T��v��C'�J�*�Z�Uʘ�y�-�(c�� ��Ȗ��Ȇ�V-�54jmJh�6�S�:y�`��bb�����x�%3YI"�!4�2sxC�IEf��&$ۈ��?��-�c����\�
n�)	|u��ǩX�H��R�D�ڷ-��Jw+8�GB�I�	$���#�jP6wI5�g�zOS�����"b���!ɤ�,��DѨ�ޚT�SC���<��a�MY���kW �`w4$�CW5�xh�XmNR+�II#i]��M�jS����	|5R���(�fJ)$@��r�y�4,������oI�#P5Hb	4��BM�M�+�J�Bb���&������dI'��6Ƀ��uur�͖���?
�E\��)U%h�D�A(��(��l�&
vT�s6�"e���'-�l�/���m��!�Qi�gӎNh��n�6���	QE4_Z�C�cZ���yd�Ѯ!�ùI���4��y#`�qHF��T��*.�N�<���q��pM��9��0l	�@�	H�/R�i9�Dx�>�]��ʶ*���M0kLa��B��C.����4��"O{`!��s0i��[!��u�2&ܦ�"R]�;ɦ�vM,Lu������r���Z���%T	+ e�*$�B�>�6��0G�Ǘ6�ХB�8��HM�$Z�9g~�P��Ȝ�,J΃Ϡf�Ɏ��b�3��N�w�4ޥ�ֵ~VS��ו�/���?7fp�9�F���愦�E�[7��Z��	$k���"o@�?{��i��V��r��0O~[D��~H�0��q���s�h=�]1�Fy�}t6F^Bh�a���X��_����i�"׷br���=��sai#���@DוsG_�_��T���Kd��]�I9Ǒ�g%M
��d�� �I�j�@�c��pCu�b�rkD����TZP�V sM#PEn�Gr�n�_� &�h�@F�D��M޶�l�"d��BtM�~6�=�%T�[0~?[�2=�A���~c�#��l���w�M�4 b�ٝ�G��N*v*z��=�~A�� 4?9*�p����p��8����E2\����%.y���"g�43�����&;4'�J��Z�E�DĪ��N#��0P#.�79�1s@�Z�;���s��B�Ҝ1����=m�n|�7>~s�'��+i����M��¨�F{K~"O���ȵ�d:��{X� @�#v��\H�vy�?{�v>?k�嵶��|jo��-�kjަ[�+�8�yI�"S�M����'&�t���Ȩl�ڧ:��C��i ;��F����fZ �ަ�e5!!Y�>M;ĉ���i�	�J&|x���@D�ZٌT��9=�1����q��ࡕH��D�A$K�.TйR$.�]��2y�̥B�]D�y��W#�T(�@�'{\(P&�tR�L�r�x��qAt�m+��� �[�V�j59��@RyC��A��P�l��8��R�!�|~D�O0p-�\㩣�%�T�d�z�����Ht*(R��±5`�t���d�d����dLw����m{dMH�~���s7y;5W�`f*�>*z����'#;��@y�w+�R*�ש��@tx��ڍ��n����N��;.~���~LIA��%E.U~"�?�?hPT�6�!0���cz'����e��59k��~6޶H�%Mj�`��كT�lۚƆ ���`�A ��IZb��
*��[CT�8����	=�m��G3s{~*0���NON#PF�N[\��� [#(��>��4]�"l��KS�$i�����7A���Z@�ڽW=O�	�=�������^�G >.Z�J�}A�c�L�y���2�qa��E�z�}L7M���ӅSߎ6.�؞�u2)�+�E��/�iG[�4�j�P�s�
�� gʇ�	m���@�H��ԁ��A�1Trh<�2|�h�W;��j�\���D�k��D��#?M<���eݟ�mI�n�	��Ի�B&���m<ͦ�zs=@�{/D�2��y1�[}=~e8�����@ӽ�p��dv��˛��s���mbH�M	�
HӡI�l��#�ʌ��<��(4'}l��{�O�ψ������[Ҧ��u��9��Pj��-raC�$�n�M���i��zcjD��lz�#JJA�J��M�<��S� -ת�ub|(9�H|�w$GM�kZ��59��~�t;��D���)�M4��"ڑ�}�HKP��1�4`&S���r#+$����ۧ����7�BIꑯ�#{��~y6J
�S����I<1۰�{e��?_��nof
i���6c�NMPf�`�h�@ xT`e�؃F�K���G�{@RzP�s��$�˅2ѥ���,h�9T_=@���
rG\]rsOv����Ȭٱ�D�ʘyH狭�2�����g���49f�����-n����K8��9��Oh�Ȍ���T�q� R I�J�풣w��ٗds��QK�s��͗�>si�����sI#�[��O�4'O�]2`��M/��!O"�@񁉵Y)[�♈3|�פ��Ԍ�5skċ���<��Kg��-������l��.l>�0[��;ڧ�{���к�DNu��"�a�y>��ߞ����������l5[%ݟ�P�� Ĩ�к�(�Cg��A.Ar\��v�h�2y�̢�Q.�h@ʤ.a�V�A���K80��s��2��2e0Lw]\2e�/��Eh�>+}Dy=��S-�z> ����뛙n)A�$	8w��rT1��$�S�rT��n�PS�l??:4ȓ@/W6��<�H���w�HR��d�H��#Y=��<�D��&���M�A���hWۗYX��	7�3����ID���%�Ȥ�Rkb��ܫA���iqVD�sjܺ͡%c|5Y�	5�	�rĬv7k�Ě�6��H�1=MF�n�r�� �"T 0�l�".��!f��WT��u	��<� ��y����;6�� 4��*wB9Q��ٹ�c���L!��>R8��K���AZh��<�8��!�	4&k[%g�|Hxy0Qam�ZZbX�I�>rT�}~�e��l4b��g��Dt�(�G��'A-�PyZoˊ�c�m��99b����	�S/��#[/���Bi��Sw�9�	��NL}����[,�e�E�Se46�6�ޭ:���	��hY+O�Ӓ��D
A�Ne�Z�!E����y�.)U�𥷺�V��9���,f{K��g+� e�,f�~B{=2n�O ��^f�@|�_�\ҥn��eu�=��?��ػu�b6�� �_�=��'�sw'�@�Ԉt`H��Pm��ҶIkeI�^��-��A�b{LSكّ$��bG5+z�ۦ���#CMˮ��-vi�7 � PN(]��}�1Pg�M9�lW�SC|$�&�����hS=Aɷyv��	�"ޘ;&�
	����L��'����M�u�׵ԍ<č2�l�z�"#{2F��s@aP'�D�E@'�&���G��V���`�L1�bH�$��K�K�"}}#v}(vZ	���䫀"J���dH�m�b(�G�{@�$G"<���M
����m��0T��,3�1�u�@ȣ�N*T�;("b�ǚ��A*%��?G[�|�	��q�e��_��?#�2������r ��Q��4V%D��B#���8q���*�AR+,\��ʬ����e��$��6�ځke�
r�����,2%������	�M@�`P#�i��!����9�Z��(L}R/�)�rq���j���F�zW��㼐�Db)5�M�5�jw���=J�]Nn��M�$:5�	'Bc�H�ڒ<F�D5Y#F����M@��Y����F�i�e��{_�>�Fϔ�!M����e�`�1��yC'���Xy.B��Cf͖1�"b��-v�h�3̞ev��uR�B*�Pf�Z+k�xc�u�0�C���e���l�H�U}oJ�#i8��#S��7���5ޱ4����喼�v6�Mc���ۙ����4�p#��i�\�ēʝ�7P��&�ǔ�ղ�B5NSt6�"�-�w'���$j�j�4��JW��x)8��rփH@��j�	7�v�!��d"5�EcBL�WI�,I����t%�N�傐�ܦ�k7��<�)L_�\�6�Lڕ�uq�"I�2��BO��L����Vq53c�\)/��fCoT��rD
LH�J���k||�6�j�C&;5]�jGh��S�]
B���p�,��Er&��R��AR*6W*D�R*�Q"8����P������a�_��'�W��R���q��{70J���zy�2�DE�Q�g��L�YP&5�)h&�YNdm�3���~|n"oI�js|��}w����'�5K��~敪��P� Z�.��y���n�J�v}?v(n�[~8�`޽Z���i���mp�`��A�kv�f�����0"&&�Kv�w����V�y#u��_�9V%Ԅwe���5�0{A�P�-��KeOiJ�˵\�;@�?*<����.��ݞ�qIa�L�P��1ʚ�\��tFV�����Fg�ٛC��A�ۮ�f�h�OL�'���rt	�$��5_i��k�0J������O.������8�8�L��8�(cL3Bz:�ǈ� ;ʓ��i�!��u�粤k`3`���eKls=9si�*j����/m�dm��zP��0Q��#�s�����ʍ߯����C�i�i�d�w=��=�(�j��M$�Y�0��H�I����-��*�n���/�#u�M�tsI4=���G�����{Gp6-�$On���*l�\�2�<�H�\uȹ�aշ!&�s����9�;A�tr�ᅢ��%T�h2�8y<���T檸R��0�YpG�Jx�����<*�U�h�ꟑ"Ge.���#/��"JR��3�iW?*��h�B� ��Cf͛,\�V��ڀ 	�k���x�R�4<��".�e
�R;B"뫶�PХr�]T��H��h\(�p¬�POj��	��H���ݚnu��Qع�(cw#t�!�b�_��"���4
>~J�)��PGT� �~����m0��5K-y�d�DL%�S����a����I5����Y��dây�(i��MDf#Hٴ�� w�70r {z�0���By���	�)�����TVkC=I*���i����Hy��a���+��"2��)�G8���CT���A,ٲ�1�X�Z�v�h�j��PEAZ�v����<��\}PƁN���tZ%�2�JQ�L��GO(n�[�j�j�,��E�zH�OX�J�y9J֓&ԞP�1	7�#�9`��#�"h�ȦD�Z��SLI�7_����iĚD��ĵ+��Wl��d����X��ecb�v_BR��u����6Ԯ$ڷ-x]&<mS7HDi"���F��N�zSq)�J99�x�Q�z`�Z�mI�������Mo����f����M~Rp�Vm��jee��֩��ZW����L�)B!X��6>I9Du����M`C,�&Һ��%7�����[-p�LՑ�ВmI���3����ˆ�*Td���T�+A�U4.h<��rTK����v��p�H#�P>i�G��#J��DֽH�S���'���ߚ������H�4L��w5\#���{j��ޔ$HDa�l5��Аc��~�'�6���d�U���)���6ꀑM�:\�=+u�ke�@�Se�M2���F����5�����]���|<��(�>���Ӛ�(��3�"�D��"��P��L �٢���eج�iyJ�,�eN��(�bm�hD�;��À��f��bm��	���̴"�\eR��da8�V��ʬ�J�]��䨫��O~����WԩC44���ꡊ�=��[�!h�1����@mYS�q���c�j�4�8���'Z2��(O�_��?'�&[��ﯤm72��A�����n�n��OG|��`�����M&���T�4Ų�hU�D�7$^�W9j;�����fe�\�L���!�\��z������&�XKR)M�v��ګ
g��BU�vZ�xy=�N`��LGi�)�;LZh�P(S�A(�)� o��*Nh��`(-�T�0��nh���H�����.��r�Љ�d�e("� �@%N\�j A�/.�x�dM�.�CCU8��2�H�
a�vGa�v4#�Dx2%Oȑ#��3�-��F^�"��tS�,�� ��ʑ"\�ٳf��\��]��5�!\��ǚDqr"���u֊#(�UCB�TG��.Ш�惇��(� )���5K�� �����۲aQ�"�m�?>l7P{=K8�vs$78|�����- 0X,��d�S`��I=�>�#o����A5��ɆLn�RK��#�m�F�;��%!�Y�*&��ִ�4ڜn�]���N������9�x�AH$��{s_� "A��D�P{(-8�l�]�V����(�B���#��O?%\]��Q0�<�&��*D�rCf�&X��h���v�Ub��X���%D�a�@�{J1ٲTn�y?-�#��=�N=��d��5=Z�Kj5�J��'�4�M�%����'Y�:t<�G8�.�6@�!A�����4�׋"j���5?_�O�CU����Bx�Z�t��h���穨�H���b��O_&���-"@�);�$n��yR�<��:��xI�t��D֑�כ�&��zn@wt5��Oe́'�jOkDM�ꐖ�k�-�MHiS7�5)���n�!Me�j�NV��A��S(�#Y�Mmڙ-J�I�S$�|�ǀ�Ox�� �A">�"m*��������4�
�D���Z�D�	5�q洤�R,��ji�D�����៑��dc�;������`��^�%D]����,<�$�f�U��?Pi�''(;svP}T`��6F��l �y��GV$"c|�+�B!"�
P�aYb:u���gi"r8���x̛H7�P6�������v~�L{�
\�vvF�?ND|Z�_�j�h�]�M�'��i���j���H��)J�++`�*��e ��^�8H�DD��5/��ʆ�cƃkT���\�"rj��O�˟�t,�do�9���ڶځۯ�$���������'���O�Df�3���X��B��hz�x29�4�m1��%˗W2�
���S�r���/������s*�c!/{j��i��mٔq��&�&�O2(m0`�p����[)΁6���4������5���� �{���a@u�n�(s(P~*PLo@�,��iP}<)�ȧӇ�m���iy��t�4���k����Lsv<~H�[t*R��Je��s�ʠ�z�m��*]0�s�0���F���U�x�O;nc���¸'V|2�J�~�kI�Oˮ"}�n�?8�$�~֑_�SS�dNÓ��!/���46F;�̵_�'�<�2�9��0aRht��~�Z���q+���ٚ!� �*����hW%A(Ƅ�k�0��P�e�9�G���恌@�Ѫ�P3\14,h�
\��U���R�8�*&.B͛,h\xa��2�B��Q.�U��_�
2\��H�D�M�h.���|�`@P�PE��{G��<��[J(���+��T��B�&G.������ '-�N[Te-��w1B� ��*���s2�:��le���s?[����T����`j��d !�����ֵ�<�N<|�~F�)⑤�J�&4�W@4**lI�Md��V����I;	'���#c'���E�刔�n]s�4���z��6W�T�AԑX��F����QӔ%ˀOi�!8��%�a�(hmA*%Ǖ"h\��Q1�X��X��h�Z�v��TK�l�
\]����g��N\L�y�k�Zd@�doV��ލI�f�lܑځ���F��5^�mU���vRR/V�ؒ+)T�5���67�'�ZWX��k"���ښ��sx<ך��r��1�KH��wR���,��v��"H<��M��J�ՉINim�ǀ�4��č��46��D�Y`H�&=J��0;�j�5RD"4�]HNH7Ĵ�d$�)��+���)4���ҞF�n��KREf���KH��͹BH�ވ�Ƅ��SqJ����rZ�۷0\Q>f���^-L*�d0�69e08��í�".4��&�:�b[n�X#f���
�e�h��oHJR%!��4w_���[8�*�{Ns}Nr����n|&DP�l�ۯ��>��{s �0��`�lL��e�����ЎЃ�x��t����� q�R�����df#Sa�o�EE#�V�EnM2j���mj�IɆ��9��j�_�(�-�k[y��4Z�E����4˖�"�*i�Lr�h?rA@�M׵� @����}LY�i�}>T�{���%-N�l�n� n�*s ||t8Z�K��l�_�n�5R��j��Ԥ�2r��.�Yy�@���4'�A���3?~d�E̶^��1����UCJ�8��S����UE��\c�<�*��ÑB���T��A�8�t
$M�H1Rt�*xm��wzѩ�&��<�~�F�l���O�#ty櫛�al��1Cbf�D��+��Fۣ��O�D�\�9q�U��n�eP#�_R��?6CL�����W�Z.i�A-�A���1wT�$�r5#_T�ʏ��L���d�zS�3)�����.|2��A�Dq�	h�	&�Z&	b~�@�2Z�Phh*{l��Ni#䣯���5A��iM�����x�V���vD�����T��tRx��pF�a��������U7R�j�hn��~��=�v9=<S��������3��m�K�݋�XrxQ䡚?*2���<`�>�Ô�\�b�C..����+��Dy�Z+lٲ�(*Ef����\ePǴv���j�%EB01pϯ�42�(��*y@�������O2 U	�����m�X�UV�FRٲxa�@�*2r��������.<��q��H�I�Z��#�? 2��1�<���������t{B`!#ȑ�X��䲃Rh��RM�3�����N��"N$rw� P|@h)��Oju����6�:']����iB9!S��y��z�� �\�\�6@�d�ke��m��e���*.e䪌�hy��A*$��1��#�A*+C+�44Z�TйSB�ʘ�u�"Р�P��4'�GK]<(�`ݪ�&`H�4���$e٪�-y���&�:^��f���U~~6mpMf����Z����lu�V���~4+vԞ�p�c��	�:�\T���HLMA��Z"H<��Գx�%h~LR�T�d���۽[Һ��;�K��̔Z<Vw���q��$By6��Z�h�4�
��ZEGWOB@"�#�] �B%k��T�&�M�]�ڕϝ�'"&�����I�V��P�&��o�b�rBqM����mMhՈ]�<wD ��Lo/���i-�@�L6$�΢9�x�F��0��)��$່ho��dm�Ҳ5$tvj��N�q%��r8jT�e�Q�L�2 c�MlS�:��r6hOhh2���L�OO}1���T"��7J�&P���C��e��O}PX�Ӕ�+M���Ji$bNF$a&�c��PJH][��4��򦈑D�f�����}X�t��t���L{�
l���
����&�z{Z����5:�sRQ��u�sL�C%�2]1�쩲��}�\y�a���\�
*N`�{]K������&�SUH@��2Fӷ@C"��цT�<�`U���(E.A�QRHy�YM,W�Fؤ��
�� 
���\
�WSĈ���c��T'�J���l�Wm��"Dc(R=[R'a�z���r��B%9�BȪ<��NI�>.�v<�����)��c��M�"���+A��&��`�1�`�rS��G1/�:
6C.?{{L�l�L}z�F	���d�F�n�Ϡ"����T3����*�U@�ږ���֍��\�)�܊��b�8mԳt�Ӂ�G�`Ԓ$��3���������g���s����]ȉ9������]B��J�)w�)�
���\̱�t6����4�S�A1s�Evr�R����@�/���hh~T�vOk�V��#(�T�b���"2���>�>�X��A�K��\]r��E]A��41�%8xS�8�B��2�1�e,Оp`!U��U
}~T]�����dݺd1t��PР���%D�ʡN�o�f@
\]+��L��{��E�9hD�aÁ�ؕT���0�Ìc�8e*QC�2����s}F�O-�;��-��]� v8��dS�D� J�����3䣪��03p�M��&�2�r���"��	�����OS�"I�L&�V.
ca�ڷ�gE�w��A��P��C#�*?p<���Aݯ5���9�ANv�U )+�� 0�%cB�=��2�����	Q"8���J�q�H%D��Uh�Z�U�.<���ʕ4 ��G�y�G�\����*hArTK�*D���3�a���0F�T�%��kH)��D%q$k��5	$�8���@�o�JUጰp��-j�$Yn�����"�:'ҥ�5���ls*I=�W���%%!�du$KyZhִ�4t�c��M֛���"K4.�6��D�C���'�pQ��ДcU��В4���1R�$�18�*ek�j�[F���RĜ�)-U�@�x�&����hY4/�T�ƴ�������H�T�iI @�)��"95("�T��m\��M��3�g"�C����:h��o�h����7O�.~���p SǬapOh�n�Y�SD���s ��Q��tIZT�P���L�.1��'7��FOaA��l`!�4*�`"���$PmX��G�zƘ��@'-l )�+�-�tM*G5�J����nCU:z��($�[5��e73S�˼���c|<�,�E;�F��,Q�i@�b�bt.nѪ
��T�j��4<����X�-�L�����L�)�� �T�櫐���B����Dm�-���7�F��������뚤�Fo�n�O�=��]�4w���UR�N�I��R1#\ h����Y�ϧ͆��U*p��"�?QW(*:8�p;�����ت-��@�O}�r\������83[(��q"��^ �6�'��'&�I(�f�r] CӁP�F�J�~�)��s�˒:�	O�^��5�ѥLi&$�Mza��TףX�0sR#m�մ�ȫu�(�uA�OX�����GRD㠚���s������Y(}Nl�����WO9��H�h�1BG�í;Ef��j��-�D�o���`s:r�r��y���)��G`�I�ckp�(��<V�į�R�h@�@.�]�Xq�+�xd ��S�<�e����u3@2��+]ED]pe�^˙ eP�SڭVzĬbV����5�*�"<]RQ�4Qb�*8�Q�J�"Tq�P�k�40ᔠ�=���?? �c�4-�FĨ�Sݝ���7e;CJ��`��S����%q���%D)����'�8PÅ�ߓ��)ɍ1��4#��]CEDd����Ȍ��"vON.��dɟf��s��庀��A�6�-+��I��4R�eu�E٢�]m��Mm�W�%Kh�oʚ`/��7]�۩H4ۮH�F����R"�yi�B4��S�e�vv�{2�LJ��v$OI;�ޣh�e����[����9>��=h]hU\�͌Dи�����G�<]��ʤG�A���.\�#� ��*������C]A�f��������J��C�#@;'�.�;���zS���W cC����S��������I�?7c���'��B��m4`6�"z��n�R{U������m�&�	I���NR�Z�ů��5����L�>�W���o�m�Ĭl44���h�6�-�5"�x�ƅ�P�1=MD��xV4:��D�'���+��B`��~�&6���D�5�J%k�5����1�K"ɰ�"Z�)�̓ 2 6��T��~��eR:z ɍ�k|�&�I�$k��|T�)�FӸ\�hq)Ri�#֔URQ��W�25 1��5)��%��>��\1m�8��������s'�G}~b��KN[}8�p�s����~@]��#(����4�O�� di�h�dV�y�B��U 䍑�N�&ɬ�B|&k)�)���bP�d;0�6"FX�_MNJr3sJĲ�S7�����18-�x�s�^���i�߃�*O{.��1��1���s}7i�F�K^D�ɎA���4��� �9i��[G�}�h�.�����1���q� �e��l��)��:�n�	�\���_�)đ>���gr<��@G2�ȧg���3CU\�
�]��k�ߌ�GJ�VA�����Y�K�����(���l�^�q�\Wc��������]�� �T	Ѧ���}=]���j�' 2�{0p� �����5�#&�
��%!l�b���=q�1��zn���-�l7�ʄӅ4��D�ҥ�4l�(��t�m����A6f�� E�&��t�z&�|И*�.�~sI	��"~�O#'���m�����0����#�
s��ey8 �u���g��*\�H*��iC2��������" �{Gc��dl�1��22�cT��R;Ev��CD]r��-�X�b���h2���4TG���*�
+���*
�"\�G���(���
%�%8y*T��"AAIZ<����BW�5U��r8!O���9��2�����9�<���:TGWA'>��(Z<��
*W�M� �O���<(���(hk�T��\],��Щ˽�4F49��n��7�7��櫝q=�$�U�uV?"hi�G"O}_�O�]�Zb��c����7A%��>[ro��?8�(T�?�(�[�d�aѽ26�>kZ҆���w����S��"@`�ʉ
ơұ���_���PrG7L}*7n~�!Cq*#�P<�D�"\yS�s�Q���40�:T�"<��ʥG*8�rTK��Dy�Q.J�͛61��Dйq�K�=r&.Kb�u��Щ(��h�Z���|:��*˂r>#$X�.��8)�~P�l5Wפּj;�k�L�0M��-Gv>@ːe����r4��H5S�
D�SSt��<��V%f��Ĵ��:���D�-y [&��kxD$ר5^����,���r�-���Aw{^O1�EcB��dK[*y;	=�F�'��s7<��p�t���+��CjB[��&�gp�xڐ��u���BH���cd��8�6�kJ�%�#սNn�#@�Ge�M�%��mW��5�<�Z���VnVFк�`�se�-k�`҄�z��7�6ki퓡��<[\�u��f��A��=�"]PdqKo`�>��k�	PPOs8Ѐ ��%��CBTEED)�������@����O�'�$-�5F)���	��#j����<�"s1:$Nu��i|u2<aI�o@�R���Tj޷�k���������P3w&��!��3�Bi�bg��no�ն��խRJE5!M�0z��&9=��9�6C&;@4Ne�H��{2�TSDR��B��O_�.nmU G��i�������[�mU�4�`v�< ��%�c*��hG} 0��H��j�Z,�+�'��QO#�vPs �
�	��Ӂ>�'�GJ����P��DF��a�F�"}�L��ET.n�=�$���9�c���PZ�o[�8H�t&��Ҥ�ˎ
j��e�Ӂ/ψ��M�������?#S)��ʆ�3�2ˠb��� ��0w���ٓ��r�e����Mش�H�7l���f��$�Z�8�M*��s���9�$i�v��Co�ķ{Z�1>�4Җ�T&	��GI&4�H�Z�P({2&�vDМ�SM��2#�˧�ڬ�sU��~Ty�)��3�A�1ͦP��s�� eP�K��DeU�X�b�FQ.J�v��rTTp���PA��Z*���.01tG��A��41�%D�*$G�A��U��V�Ce��tAJ\��CJ��Q qu
8!H%D�0���44(�.��8��B�Sdݺ)��ʬ�\p�ۓ�p<0�e�~pPʤLh]T�Q��_��̠��ZY@� �" \Bc��Q�^�?o��e�[/9�y��U@�L{&�H��G�� ���"i�&�:~��"!��6����H��h&��%1�j�}z���	���3�j�&F1�|�w��E���^�(,��BSv��R$�c�5�?Q�R��BЊ�
&.<��l��T�a�"<��ʦ�*��h2�Q�ʎ.\�䨗J��Ɓ�ң�2�(` =�{A���#��Ў�\+3��g���Y|��Œ[rN	-LT�i�ċ�Q�����pE���zy��B;f��]��m1�7h���n	<M@�x܍b�-y&�F"�ŦI�9d��ט,@'��vl��7�m�C�i��e���y�ڑ�m)��q7��mbLF��f m�����oJBk���0��mH&$�j�����{L"M=T�#�%8���S��[�I�D�"z�[�$u�ӡ���6��CL����I��ԍiL�b�΂"��AY�+=�H�K�4��|���$M���ұ-��j_���v�l�AR��C�#���ݘ0�c@ŷ�ꁃts�B;A�I_\��;{O[rp:�MT� ��a����h�EJ��hU�ؙ��e��j��f1r�j�m�J�
�0U�qrDģ��Sb~��K6��ͧOW����W)@��4EJͫ�md$¥e8�a"����V�t��$H�F��5M��Ef�D�+�A��7��ÚكM�$D�7���ˢ8�)������@�{�s����S�⒰�NA��-���OC��r~�D��+���̜EhE\Á����"\��L���x`!J��WQ]ha��kb��UX]P��sU���B��h8�(���N@���S����^Ҡ���$mV-�<�v<ж]���StL���~��7D��X���TH�D� P_�ͭ�\�̺��	S�%L}<`���$N:�ӭ����C�JHLj�_�N���&�;fOΈ҃���#r"{|@�)5W�#��J�O��D<���O��]�%7 �$ݾ��F	��L}n���7��n�t7Pv�
����"n��`(�!K<��r���qȻC�T@Nk��A�=��Be��
v�Q�G.2��E��j�AP�M�	F4*8��W4W4P]b*#� ��G�2(�g��ϯǋ�P������ ��U��k�U�Р���*T���c�8e�����P��T��^�]��������Dqu�c�;`������\�YD��P _��2���t���$�H��"<0ʣ)m
��2��	@
��. D�P׸��t�v��f�2�ցH�e�1=�Rp�qs�Nt��`�k^�p�M�AR�998��I<j�L��`��#�"�yթ�'��v����ᷪU�>�
>j�>L`~���8�CMb�[z�#��7n�l-�"�B��Љʐ<�)s��}~h2���C�Tqrb����\�eQ��U*8�rTH� ��UC4.pR9p�� G �)���!�A4IN�kI�"Y��MS�jcI	�Y��p�Ȳp5��%�L�m4�n�N0y&���H�m�> kϑ�zWb3�e���9�N=��G?<�p�*u*p�⩕�u��Kbi^ڴ����"jE5;կ)8P�뀲� M;7H4�
����4����6q̵���4��At�Ȗ~6myJ�y9j�4��哳jBH�J�#HI�:��JCIH��"t-�5H�'�Jv�C��׈�bjs��I�&���W��ٗf�e2 4�jM;7J������Hڛ�;�ǖM�דr�V���>zø����_��2!�����gK�J`D&K&=��lm������C�$.�	�m�Њ���b�u=ɲ�����cB;���`ɍ֛e��ON*-l(9%<�ؠ�Ҍ<d1pI�M��
�tz�G"oT�bf�T
 |�.`�P:$��*v�MHj�[��Bc۲4��>��K�&9�[�3���u�X��@	
�尒���-i�(LA�;am����(00$#vLi���
��H�ѥM����A�u91`�$-8�*�����8S��Q��heu�
�\��K�����=u�a���Hש�-�[2�����P�y��?h~\���s}<����*������ r{2�B:S  1S��H窴T4 ^�hGKK�Bt�rx��y1�r=��R��PG���)ѧ��^���݌� �4S*�r�Պ�D�w �;.tʟ\��eg5<�@��Y�����&KoW�O�T�>74��� ��\탐W=���?'@ҒĞ�CT��5
)���O�m��Tr�e 3��"yL�L�'%˓�0{�"7~8�rTF�pm8���H�}�i��As�� "���#�{hi�&'��݋Vߓ�9���҂8�b��"2��Ț1r*D��u
G.�Ȥ�	P<q㈕b��H��P]Tqr#� ���Q.Дa��QWPhbDyG�A��U���PhchQ.@�V����1�c:
�.8z�E\]�qv��v����~2\ ��0�Ԣ�#�)���A�V��W ƅ��
2���\�;�g&�z�)hhl�"2��\0��(k�E~s�~٣���K�hn�>�Z��Ԫj�%��X���� �.ǟ�Zmt��7C�D�u9jh���9`�i��<��'8I�'�nSM8�Mj�$�����0*:@ �|�S�� ӑ�����1�f��E9�^�4����^`�y&=Fݍ�'R��es<�񔧌�.(``@�8��T�*$�C\�*%G4Tx�A��
�.Dyhc ��J��4<x�ƃ%��J0 �	������@3�|ڃ[R�����CU�1f�H�[�E��TΥ��:�`Q���cZ�^���Ԍa�z�j`�i�hH�� 8~56#�sx�6���[������Q�2�2��������!�H�[�&��K"� �ޔ���T�5�U�jL:9�:����^~@׊i�E�)ԃU�ě8�2�7w�RF���ۉ5�!㠉�w+�
ja7�e��y�:�l�T�宆���&�"_�Ѫr�Ty�F�J�"���֐�����j�em��M(�Ƕ�5��[L0z��KpIjL+��FԤ6�6�ͤ��� �9&��Z�$�<<�l���v)��)==�R:#�K���f����8dQģ2�\�A���=�n���9��� �(e��R�G.\PǷ'`�Ϩ%<�����Dem�����@�PZ19�P �3�LҲ���wa&�Ƙc���2���ױ�C��I!jd��ajaC|� 6�й5�ݧ]� ���m1�`D&�l�S���7fʃ�!NO��hDd�wg�I�ϭ���3v�U�<e I��m72��8��Z�� .�� 2{���� ]���8���"����ʜ��ꧫ�*G(�b�45S =�9�1V�e�6�ʚ"\�ī��<]��#���Y�ʀb9�#�D�x�$u�d�0�$x��J�X\��)��m(ƫ���;4E"`���E�{=/�� �$~&گ�7^�<p��c
BI�Dkd��+�����M_�����zc�{���:~�0l��'. rs�U1d<�w5���{B`�p�9�jٛ���&�I�|�j�-�SJBw�IF�ө�kJ�G\�Bs�H����AЀ�$P�4�A(L �l��2�1�P$G��$�[z� [��&#��v*s� yl��ٖ��:`��b��ߏ�l?@.D�e�(��8(b&��X�r�˕"A���"A��E���+�Dq�
�	PTy��W.�J����WhhhhhhPhbA��41���G�\�hl�\��c=�&PМ]�� g0��<��A��/�����P�{G8�f������а�P<��
���J�]ʕJxa�6P<�q� PLl�Z���e�ɍ5��a�9ͪDT&$6q��(�1�:�-�5�B���*�몴T�E"8�|�$&��%<n�x��b,��%�8�(���ں��0�!�W%+���qRib	�Ow���(�R�"2b"4�֚Hy��:D5:�-��ж� v# P�v7�P�"Dd�RL�A���b�h2��WPhb������ArTMU.�x�B���A���.TqA�MU2Д�ĦL�.���w���fUNl�/�G[�����jčbN:�ǩ���`�v0X�	T΍�3h�H�H��M��H�,��5��V6�����V��W���&ę�SX>໩�+�Ʈ%�r�I�Q�Ą�oI�5�Mj�z�S�%ϝ�2�LH�H֦;�)�f�26��NN-S����A��Kah.]1~�n�Y�G���j�IV�ӠH��S(S����q�j6ޓ$�"ȚT�;��[�i���`���):��$�0��֘�T�c��.�Y[��C�d���6��>�#������Ť�v}J�q��F�I�2��ebڔ�Ѡs(��٨��HHI)����h�
#�"T��<�rSȚ"\����� �(R9��0�Ç�E�nN�K�2�]LJp�8��*D�SAs*��F���	1)t���dBm��F�@�a٪rGh������'��ԓ��`���9�A.�b��0��E���to��N��0��*?\�f���nc���O�j�\(0c�s}j��-�[� ���j�_T�	�M��H�|��|��j��el�Р1���L���� 1�ьhhs~�EU�T�1Pd��QhhR�<��E	����i�Z�\��D�3�h@ᖃ��(�V#�h}��\�4=�D�p���s��%�_�-�����Eoj��Wh�#�h}9�3G����q=�m����+h�{#i�SCc�v��.�<�j�Ii$�~���n�]S��q��;j�>*�D�<Pb&�@T'$���6��a&�sw4��fK^�H�F'y�Ќ�ɫo�ć�p�֢��P.<�N\�p�k����{��6�+Tsw4i��]���1��1l��|�*T

��'��{U�n��K�_�9�������"��'�}-N�/��R�}Nr�g0b�.\��h2��ʥʘ�*%փȐE\��N*�p3�p�~.�(�%�K��PEA�X��X��X�TQ.�]D�CCE��\��H�*T�R��R�5� ���a�pB���GJ��*.иʤG^��Q��GJ\ �Iϣ��l�yU�4.On��
d`�IZ,�D��ʫ�sPNt)�R���� Knnj	��`���s�ɔS+��T��j���UQfP���D�#k�N�MR�	͇��]���&֤��I��"���W,����3�rxԖ�X7��i�Ē)�i�m�;��*0hj�ڮ�	� :�~;l�($��I
�(
n�QfOZ1�r�ʕ%hT��q�H� �%�K��Q.�]D��u����S"JqQq�Q�Ge��P��� �����	�S�9��Ѥ�O$�|��e�Q������X57���|SnG��p�|No���	$�Ց�j�~�~i�r#��N7I��e!����Ȭ�Md���j6ַ-U9H��+��HM��X��'(��^vx,��2zLq	/��L�oBN�-�S��򳈵b"0S���ҥZ�T�F&�H� m[��M"b5�N�da#j�o�K�IXFޚ�5+���$k�DI�`��9���5�eBjr��֓I���5�L��:��ۤ�뀲h"p���c|M5�:"I�b��WRT咺h�ܑ8$i#��')����[4���̂lN �~X�ѢA�
��2kL��*;�TJ��a���Pvs[��\�p�A�G�8	�2z������)j� �蒴%G.�+C �S �+B�*�~�j����		
l( 4�ɓ��H';*7i�F�m��I`�0`H�����4ӄ�O%NNs�����U��T���IN���Y(""Tx��J�P]b�"��}R�"D�)���b�4�oZӠ���!�����#^��G8��̠�v��%D���]B��i�VN������������t��d�Qh�41)�J�.���V�\ʤK�*Tйr�IO"Jy�r{.��]D ��
��P}~n��[{b9�Fy�����L�!/n��	@q�vQQ\��P$� 	�S�-��щ#r!����#���\���6�}?~l(vD��7`� ���r9���6�w��w"��V�i|S/����A� �V2�u��lQC����y����[��@�h¤a���O�
�n�ï�M�a-9�����4�)��n�;.GL~2���Av�����}d�㒡M�(��Z�"vJ�<e8e�s��u��j�7E��O//����
�f�h\��#�.�x�B�����D��1+�'�g��`�<��%ʘ�S*b%�K��PEAr�.T�ʘ�S*b�L\���1� ���C.A�"D�#Ǐ4441rk��1**�#��#�A**�#���a�T���=�(��%Dy)���h�AQ��TpP�5���J�\�����9����D���aVl�G.0f%U2�R�ٗ0���[+v�@���-�����}.�`�������#v���l�¦�Ud�<|�����ڑ�ݒ�-l&��ŉ��p8ͦ�CQeb����Z|ty*"O�4Z��c �9��5Zw�s*V�)UP�1��b��.B��(�Q.�]D��u�%�K�B�*�Lh<�)�FK��q���u��#�T�)S������~.)��;�[�j�L($y�,Zg��U9XLx���F�,��k�C��n<޵HK��9�ޓ��g��5��@�~$0ktM$�R�����S�.F�4-���m�ͺ���DCƣZ��0Dmzp�e)���H0�4n�	���ש5�;<[кM�SH��C�L�J&�lF=53�驞é��Ác�+����&?5��	�f�;8G����yMf�6��A��]��&�4��&���.Z�,��)��|KR��*e�5�-y�^F#]xY4+&��Ou������n�Z��à �ګ���)���^P�:=VD����#�S�u+���u�,�֩"X�����
xP��ZڍL�����˽�8(1��a�-�{�)��8���p�`a�J�	��x�g�C.8z͛,\� y�qĠܚ�dCbF�i@�Q��2	��l��zHmA�DD�n�4�A\�(y��mId��:�0���n`n&PPDDDF&F:D�7>?>L  $H� ���� ��"E����ɅDEbD	�S�4�&�b���zN4 yu�	Qp��@L*>X��"'�#��M&�e��oӈK���R�%<�u��*.�Ĩ���erH��!�f���r{l9�=��[T�*���VqƄ%@cD�)�-�E���a�ص9 ʎ>�<����]-ȑ�T׍�s��%t&>�H��ڮh��Y6�ѭ��S�C����`G�����|$�߄�	��W4�$H����n���NI�MK�N�uENt�'�ʒ��Ph)���b��L���	��ە�pQ�8�����4r5��j}=t6��a�d�.sUK���G������c7#�T�'�����?~D�r��9�X���1mp�B�_�V�9-��{e�PhcA�Eߌ�~2�a�G�A͔K�N*�pR9��Z4 �SB�M�*D�R$K�D�K�D��Z*h<�SB�ʑ.T��.A�ʦ�*�\��� �&1��b�,�F���-��<�Uq�V�Pд<1�(����U~2y*��
�� ��(*D�p�
��.<�)s��N�j	�Q��80�8aG��	��L{Ns��nFPx28�&�kU�͔IZ(��+E�򃲧ш�K��\�����1��ֵ�l���4V�1����Y��Nd���@��ԁ1H�~$#��T0M19bH\H���N�=i�l���/ǋ�>��#*���Q.�]D��u���PEATPEAV!Ar�4D��%��`��NFb9tH��#�D��y�;�&��jڃwh8)�A�:�&|&�vl��8JvԄ�+	&�'4 n�J��g�g�n6�5�n�(o������I�L"X��$����D�\�ySz�FtNMOP#:�� 3i�NMo
"%�6�y�nH���5d4��[HT�&8
i��D�)�[�z�NNH&������7��γx�d�SZ����+R	+�	�!��ta���:��T�	"�ȦZ�;�8Q���D�;�L �7Wj�O#{j�\W�jl"R�Ί�yОׅ�K���;,J䵑5`6t�8���ƙ "�{��I4S6������?y5��jtid�׷)��58�q���`(S`���)mᖁ��
8e�0װ���#�=]�D��;���M�>�<�Wh�2���?<��q�ˌ�{r[7"z�Fޮ�DjN" +MB\�O��F��S��N�:5�(s�'C*J��m)������
q����u�ml��ܐm�$r[sh<���!D{e[6"As(~x��0`���#�~))��Nl'�hTqR�ʗ"h\�+CAs�.U�'���Te��q�<Fm%��(>�h��Y��N}J(����U̮erL����*�?[n��Pv\�C��d1�;DQ�O��eu�����:���V^1�����1�2�-{�u�j.��ml�j�>;��>���J�䍂C��#knRPl�r<�`�	��x�0�t���ij[X��j����3��y}�*�G86�h$l4��w�%#rD�vaƙ��e~�jn�����i�,�-��x�S�5�����$�Ll�\T
�U?hDH	��J�qS�DV+��Z�6Q˴�[3ɜ$M0����[.k�9����De�a�3��fJ���f�m�'%5ʑP�J��v����)�ȣ���TЃA�K�1�l���EhT�K�D�K�AD�1�X��V��Z*\�%� ��CeQ�˒�Dy�rC��4(�.G}~��]���hy��<�@��%EEA*"�.2����:We0IϩE��T�����e)s��*Dк��ʟ��
 ���H�?=���?n�6�<��	��
.Ī��Sۓ�Tr�H�<��� ?r}�h22籅�T
��ګbF4��#t��G#lӆ>�5@&Vˤ�9�Z�:�$,�ɋ��^�M���H��Y'��������:
;Ϛ Ϡ\�
F���
1q� ǀ. a䫏%\��$��4D�y���\�*�"���*�"���*��1SB��8e��s���G\����P���̪GG<�	�m9��N�m���`ۥ��$k��F�:r0tDMR�ySȴ�~l˨(/���i�Ď����H��,��rAe(c����d"'�f"rA0��`�j�5�BGt�F�3L�~VM�M�D�kF	�h]X�;�$jrbؚ�̵H(��<�;��+7�M`�+ ����NX+GVB#���'7���"H��X�ZOY	!���i;)	m���By�@�ǀ�5@�G��&��I�&�Gl�7�%�&����M�1��L,��ɋdM�h��	�ɉ�{|No	�0w��S��@j���v5Ƣ����!��d��~whl���$��jX:�[�k��hmIm��B����̓�ШR$#�  ꣋���45�<0��� KnT��.�Í�R�2�p�
}Ov� ࡈ��8�)A0�m��o��i�Qk�b�"t<��('4'9�{�C/�O6	�z��	S����`bH��[Pn�Oϋ�����ʊ]���){"ٱ�4V!�bD��P�"�"�e�PD�M��=��a�)F?#�(ࡋ�cB�d��/��Q�١Gs�HDX)���隉�s �Phe@���X]URZ�ZU"AR*-
v~< ���UG�Tq9�Se��1<�p&#���PJ�c�8�`ʑ�1r��U����u:et�9D�Gh*{<H�*G�%[p�&����7��2&�T�z=J�Q8�
!Չ �s2]@0� �9�a�yܴ��~j�-rG([~l[�j�͠m3S��@ �w��@����1��^2�m�א[a�d�$�[J\����Z扲*�d`څ��&0��<2ź��r�֋�!�vE��n������6絛�_Z4�?'���MV�u8��t#Z�y���s����z��e�U+�V�*�]hb	Q4<q��8�ߌ�.й*&�*�%D�v͖!Ar�1��6l�Tйr�H� �&Y�f�v�]����B�1�`��*T��M�GJĨ�@��E��8��QPJ���<��S��@��U�U=��P?l;(9�^� �`G��h8y���6l�h\x�[6l��m�����J�q���O%~Bƅ�.�Q��C9�'�7g�"q�� .�`�.~칲��F�j����ڭ���y��vK�&ڼ�L��#<`��X�=A�1��,��j7,����-7��˱��@�Q1�l�RI�'�8ك������2�ʦ����Tq*䧑hASB�*8��ʤPEATPEATQ.�T�MJ�)�G�.x0c/����.���E�%~0��gg��2D���v�5�$�;�Ɛk��!#T�4�;����HK-z��JA�!,��w#yRM�Il��)l��ޔ�����s��bt'��GZ�&������jNq7�3X�H��,�$"�B���5l#N���;`m��ж&�2�L_�����h8����0�HC�j��F�'	�.���1�Eu��ܛB�&��$o��n�|M$Rě�q�խ(w���j@I����I6�&���4��g�����,��ǎ�!�����G+�ԍb?+8
M�1Ԓ�[໨m�;:
jSI��t�T������6���+1�D��'-TS�"�렖`:mP>_� |�- _���bE�\��S&k�Z-Uq����\��m1N�e��˽��{G2���F2dRPϢ��߆=��8���5HȒGF�~�X�[Vԡ���~���e*����1����˯ʗ�U5m��sʑ�}v}sr~���[6A9��#HȈ�Ҝ=�*U�er��A�E�bD�Ȑ\���R�<{�젉�hm�e*9uFR��u
��
��2�͚UKǵ���d�����p1�ϯ��5��Q��#*��CCT�J�\�@�ֆ..��ꪳ+�)P�b������[C�<� c�s�A��T�4?*���
< �zО(�T�w�T庪����pURp��7r��-m]��Ck��Z>)� eI�G�����#"��SA���QNJ�D�שI�%�Lܦ�>%���WCt��r6�%z����F�"rD~))����1�����Qtȶ	u8�9jأ#'��7@9��-S)G��������9%��ZA*(}�[t4?Eh�;%J��ymr�t�6�uNP��0P��<�	��Fjr�g���;&9���8 ���he��� �����.J���U\����Gdᖅʙe�X��lٳf���&1�6lٮ�k��1LAA�1��<0���5Z%D�TK������k�0���<��(��"8���J�)s�<e*�ʘ�6X�"�?=�Dк��)R�9B0��a��.�� ��ʃ#�����[5H��#�v}J)ɗ��=�T�1s�ɕ�`��L��%7r8T�Zjp,M������<��P.Zڻ��A���0r~t	�w�9���e���N��Ȓ),ƂF��@��޻<�����;
�EUb�Sȏ4 �u!b�#� �%�K��Q.�]D��u�%�K��1SB�J�)�IN*Gdᖄ��4Dp�S��G.xaw��f�T�l��l�M�P$�`H�R7�ӳխ&��9e�y6��!I����g��7b;vy9;u<�~�yF��1&պ`��T\��MH�M	�6���"D�Y�t!�M��k����w���Ԟ�5��S�I�!-T���Z5��`D��F��hD�1��U(�jM��c�jWI���!M`t;I��!M`�T�|�v7y n�'8�Bh�l?$Yr?#R;��qȲ�� -z��CU�	�V�Nβ$�8u$N&6���.�)��Br��bX���\�ے�N ��.�#oM�rb5�Ii�zOI��[r$�<�d(X���F�j�.�n�(w�K!u㽯4ri�:E`�d�W7"�]e��T]��J��~2)�0�w`@��òۘǴtpB�>�dS��OcU]h2�`b�CD����9���=SI����iQ��Ў��AĚ[{c�w�6��6���{A�����q��o��B�Y\yS�!�����"D�K��PE�r��1V͛6l�� �r�H�"D�r�G��*D��f͚&1�r$�Q.@�s���.<���)_�)���x!�� q��\��SݚҠqu�CCT��<(�W�m5���#� �]E�e��E��x�BQ���Dy�}~A�ET)qw�(��@�*���tS69�~"s{NG �Z�ǻ��{Ԭ�}-N�\(�����5�FNo��ɧ�0�&�vF��/ѵ�q��9�0,��G��E�7��Y�׍�u���H�rT�i�[.<�\m:����Ml�@�4��m�'�jSd���i�"<:اAAR`'�w%̀�������]��L���rK9�G_��p�O{S�υQ�UNFR��\��3=��.l����444�7�%�NVo�;7Q���5�D�� x3A�G�.�\��1�r�"J�T���
�e0���2�R++�"D�K�D�1LA��X��X��X��X��ʥG.J��*D�r ��챡r����bTLJ�����������2���f͔��"h\��>�;=�Lj��Oۢ�?G.�����\�;�
T-�c=��\��t��8����a��J��J)�'�B�H�p���=̮<�3U=��#5$�����;Zk)���6%?Pځ�-{7,���M���V����dH�51)�ubP�$�	�>l�#*<FaGh�*���9U��.й*#�Wh@��$,B�TG�Dqr�L\���1r�.T�ʘ�S*b%�K��1SB�J��U�N*.0�&��"b�ʑߟ��A���E˕�ƒkjB47�Pjq�A�F`mmB�T�ܮ`mL$oL���&��A`6މ���`mkd��8����Gv-�R�TV-RF�Nڝ��c�����hV6����AȖ�H�i���j��iY�6�cP��M;8SCW��h;�f���Romi�xך�AH�'-]�Z��6	iȉX�+)D�E#��^B_:+�4�@���Ja�!H3tH��#p�^��E99~ރF�D��#��L{~l)�R�ג�'�f��4��M"tL �EN򲐦�R�	#̤ے�JQɂ��׃W�u�q5
Aj�.Ym��q7A0IH)��n�`~�W7B���M���1C��=VCSA�.k0 zҥ��TFCJ1��s��2�����rx`ʎ.8�x3��A��v~rO (TJ��G~2�\���E̗s}}-0hl'�ĀĚ�jyP�ə��.v�1�u������ )�����m��6h��DйP�ʗ?2qR��V������b�ȏ �Z-�6l��
�*hhhc�TйL�f�R$IZ,�C��->�96L�@�UUE��r{���a��T4Z�N44#�<(�W�4�*y
 GJ�0�A�K��A���.2\�q�R�T�ST0������J�ꪬJ��+!]�@�6^M2ՋU��� P�W��MN:� {j����W6C=�g�ˋ]���b�r�N*l]�� �S�$PPy��O��2��-�NS�._�d�tk��;6EGp3�
��@�Q+U�4���=��CB�F��-�Q��N�U��0	O�O=��7E9V�
[.ql���;S�E7�nM� %�RR$�M�G��}2��S��2��z�y��Kg�-w�'�6-�PF�>�(^�OG�<3�Ml3����<����1�u,Р��ʚ*Tй$H"cA�K�*h<�B�M�T�r�H*D�4LA�K�AR%ʑ ���˿8���v�Ǖ1rCg�JЩ+E��#*������h��.�2���C(hh��!hcX�d�V�Ǖ9'���ާ����PLl�&6Sۭ5���%�2�~G���0>���::���sC�������~9̻��g��D)����ePaT+�J5*�<�+M����x��^���X�(�lG0N5<����e�C�T���5e~�w��������\��(ݺ�HF�`ս����]n��Lhi�N!2���:G����'�4*cB�4Dx�A�t��TЂ��4 ��M*hASB�Q.�T�M*hA��#�WJ�b9uM�O8����i�sNhG���t'B��u�މ�҅���yH@�)���,���7�"�w!1�e�����	�6�6�^M�1�&�(k��rF��y�(_�ě�yk��<��k'�^tL�M�pە*�M�Ǒ5Jk��$����6+���.T��8	kdM��Zh��q@"��DЉ KR��O94��,����C��li���W�"�
�&�LBi"�j�7�ԉS�j�P�2�<�k����C|1<x��i#p_Z�����NX:�94��.R��&�FԄ#�ժ<wM\D�3ĩ�Vy6���ѡ�wY��i��[M�M#oM��yk���;��W�RG5�t		�+c�*;M��58	�r�� �6�_��.�pS�R��<��J�]*�*�J� �6S�� ~Dy��? .]� H�N@�h�1Q�QU\xa�FR�p��k�#�j���$ng��^��% )��RU���c̀P�(l�44X�J�*2qqĴ6Z}v���T`n��	R�J�*�!��&�G��s( ��\�0at�D�$H��,CD�&Q2��%�A2\�V!����5�&�sT���t�3�
-q�G�Ҝ]�̡��.\p��8�3����J�f�Ce�R�T��K�B�yw�%�a�\� ��P�]8�S�d.�@� \��@5����s�	a�h��k��A�`�i���	�K_e�C���W�Q"�z��y�
�sdQ�|6�%���A���?Y����ޔ6F�R�{z5y���Xa�Hܬ�+�MN����қ���wi�j�h0s @~@O11�i��K~hD�^)u��8c��u�:�]�8�G�k�2'�漎:�O8���1�Q�LBЩ��2���p�g��w�'� �\�;�\e8�8�$�O�E7^�?* ��J�.�+�-��(TЕ/�D���v.B�
�?>��}{\p��4&_���eʎ20��t��.a�*�4Q���4��4.T]��:TG �#����e�'��2\� �r��A,�
&��"b&�ǒ�YC0���THx���\P�/������} �n~Z6:�(0.���LD�(ca��������[~i�=�6''�;6TZi�(#�s?l�~CT�B��>�J����.Pg)�eEK8"�J�5[
�ߟ���ϓ��Z��h�tq֬��ʛU%�R`��o��\�Z^�[�OdG�
;
�E�Ў�����u�S4 ��#�W8���M
�y��W%<�)�G�\��.ϡ�#�{ ��� a���;>�G��`�_]�;-����8��&��#�d�:���v�S�ͺ:�~�i���Mi���8��ٰFdc'����ͥ�m{����F�_���rq��Ę<ڎ��&�����5�9�RZ��՘8Zo�h� �l���Z�t]��zz��ͻ��_M��ܼN愚��?J'�jlX�V�4BH����i��o�����1����%@Cb���6���t%��&��Ф�_��e�C���;��"&���1�S(YJ��u�!3��5�Ok[�f���&ֈ��i؍NLvj���i\�l�uh�L�MSʔ��fҡ��˱"ĤY4?ѭ��Ko� ����X���򛈀�WNoH�����ݳ���(Ց��~޻�R�&�ڠ0	��\0���`H�E%`Ì8��XЩ*8�e�3�Z�T)���-�0ᖇ��.�xS�;�!G��2���)W
n�#�Nf����̻=�a��`��8��#�h~ЎeV�.B���*ED�6Q4.<e(����t�R��x$�HPe�pR;T���9~��LD�͚& ��l�CD�4.\�����йr�1���r�.\`�B� [n��mT�2�6�x�A����Ed���C%hG{�?n��9G.�RP� 
T�1r9��� [vG{�+B��1V��#��R��*�"Tq�G�h�jv�U�l�>�9�OhJ��3D��OK[UNh���r>-oG�����z<d��l#�5���5�񻀁 FR�
r$Ll=O��Ehu<�"`ڑ�,��RrI���l����0`U94@�ސI�OnB%!�?Z	)I����\tb��m�Ԩ�q֩���H皭5͕���m�� `
�"�s��c�=��(i�ި�ӥ��Ǔ�
v�y�]2(�p���Ǩ��3h�Gc�E�Ol
<n�������$n�&�� ��Pd��A�-�J�e+���hl٠��b%ȕ4 �U4LTe)p��B�͖��2��J��Te*㇎
d1tGQh��-���������hhhK�2�rW*D��u�!Tи�V�,B�R+("b�H���D�q�Q��e�B����|�"w�;Ėک� *�������s����t�f���\��[��șh�'�8� RP��% (2s�*�%@RXƉ��+�=� �NPj�n�QUG>#���F6���k��l���Ǜ�3�������F��3v�!��!� R�R���9�?N�r�=E�c���xᖃ�Wh@��B*�W2�t�B	O"Jy��D\�@�s���%<�as�����J�(� �%\�����1���e�����e����st��T�n�=I�j`��P��{T��mc<��Wl���N~s*0o��cq��<�H��Ft$MF��A���`�&/��!#Sn<ڬ�D%a9`����r�&�)�������ZD�)��OmWA���5����DBqI��d��M��洞�&,��	"�M�i������RZ����X]XFbR���������c��BQ)���5ĥFF���;<T���hp��I�"j�m�;7�u��vLmI���� $X���ra�d��ikHJ$j���F�颚�$t'�)ǜ��3K��܎��Hִв!+򻭯6<\���$w4,J�cq���_s��!��&	�^GF��*tF�&"�٤#w�A+� ���\�r{8����Ƿ����?d��%8�r�*h@b9�x�@���.y*#��J����q�#��:���`	\��G�\�b�`��=� �Qv�ሆ�\��T4,\��&2����~�pF�g&�}	j4��EB��Z�G�[i�����;-�٢e�4LA,ٲ���#ʕT�R$Hh}0c��ءB�8�ɒ៪�@�V��@
����PvO[����*DйRV����*D�A��Ȩl� ���C%G.e��&��U*8��a��rz)�`�FX��b���
J��O\�f�ͺ�vn�0���G�>��?*�Ei���@�b�"�#S���[w�.j���C`��L ����G &�4��G�BdK!$i����PP>y6V��x�5�K%���]4x�B`t�t7�H�F����~Վ� &����T�0&��{�N�'�*�&6��3KZ�� DF�j�%j�X����a���L<��	�>?)�'J��@Q=�T)s��8�03M�3u�b�vf]@2�R̾�~l
l�[��Kg���; 0[{L}}O~{[G �}��hU<���l���Q2͚�UK�2�	�t���#�a�*�<�	QP�2�Qv���L�.�ʤ�G(S�:䨨h�42�CCCCB�eRQ��A��8��1��H�*D�yR�H�*D�yQq�Q.ALA,�\��5H�.\�$K���94�	���L�Jq��m̻��@�B� �\c���'ӏ�G3J��Nsl#��h~<���J���J��
UFA~[v��q�PA�>�$p/��i��_O�)\��Y�S'��s����(9���4��5\R����ݗ=T��B�ߒ�r���8��U�B��TK�
�Щ�
�y��hAR���D��#�%<����H�<Щ�N*�p���H� q*��2�A���00	�Ɓ��ǖ"I#P��i�)�)�-҅�P�h�����? ��#X����CQ=�+��u1L��:�D���&�!>���cf�Q��S7��QL��mA�$�������⦩hI4LYVk"�n֓ګ�IB���'$@ͧb���V;:�D��^ k�F%2�D�-D�|M5�Rz5�V2�&��D�w��I�Rս&���cHF�'$��#I�d5q:&�b�hm4/�$�Ĝ�P mH��Ԕ��B�D�6�����mx��j|�k���*�	�;���m�#���Bm �ܓ����������i1�o�I�yj��&����Չ9"j+�栒��WIJG�O'e����!,����h�D�,��� ��{vO}{{s )��( �݃-�;
v{T0�ۘ�������s�`���8e�إ�Q.�q*Q��T�TH%D����\�0��A��GJ3C�ʤ
.q�����%~��b��j�Dй�l�ٲ����bm3�œ^ޑ�UJF@H֚N�Cā��YD���A9=��0"(n�&Y��f���͔45� �%H�.A�.\�1�T�SBT�.]���б�r;�g&�{ۓ�Tr�����u����2�R&.B�4H".ePÕH�<�ࡖQ4.hyQv�E�#�T0�Q*�(f�*�v�`� .��1s6�E��#� auIC[LN{Ph�0vJ`��t6]��N.��2Fmy7�kbF�h'��T�Hֺ�E	�r%�m)�b'1�br��ܯ�N�[�1b`M^� r��n�ͨ�9$�+�O7W8���憽ٵ �*NR��&�"EL0n���"���kv�2�s~j�4��H�5[-����~��֛ʒ�.��l.l� � b�h}8)�	��<1��Ƙ�Q�c���m����f�Kg5A\�/h��� n��\3����ȃ%��O}p5�D�z�OLPTquL\��4)_�*.f���9� ���QÏ�K��0�	Q.2�q�V� ����A�=ػ�G���������a�+Q�~)�ʣ����=� p�T1�W*D��r%�1
8��� �& ��Q.A)�˕"Chhhhhh����{[r���)r�H�iZ'99��F9;O*@�V�s)_�..�ЊЉQ��_��xa��,�h]f�$�J�]Q���TT4#��rl�9����jt���<�q�s'�#��k��C4'�^��?5['��b��2�iUP�P�P$v�������.2�Q��"��Щ��8�qs-�\���%<�)�G�Jys-��?
2q*�q�^�#�~.	�S��aH��#�~.���`D&�>02���A�dj/��T�b~F�"z�^�dt@'���l�J��r�H�Z<m*z��Ԅ"kr�YZG�ݷyV�B�`�~���+6���k��$ӱ����8磆i���5�S��bYnM�&��hI�MGb4Ј�h_͏�&�+)F��ꐘ��I�W�5J�#X�V��+eI"'A�mHK Y��D#q�i��!�8կ'-V&�25dRF���y	�m�f1X��5�JW��lWT�U+|KR����I�Xj&$H��C�f�wҀI�&�.THj?F�Q�rcM֛��C�"Y���,�I�P
����h]�)�#k"s��'��&�����]咺Ħk-_��Ě��Є�k�M�Ո^RM�p�Ahj'�CV�Hb	97Gm�Nkm��e�����#�{}���� �C	���߃r[}vs{.1+�'�*��h2�Q��%D�TH%D���2ys(�D(�Ƿ�w0I@
�UJ�P��@
8+���q���ʐD�6lО2�0 C�O��I�Q'���I��96TM�ȁ�\0���JG��Rx �t�1B�6l�T�L�e��C��b!�"Tx�BT��<ƅ�L�b��
��cB�.�nbc�Ebo�Nǌ��e�&Y�*J�c����%hcB�*AR&���Uhe��C2�9�D����j�v~�b�Z 
D(���P����2��U��M�㉀b��_=����M{���(Z�M��6�7t���w�g��܁�ԍ?1��,��D��rV0M��A'�Iev�h�H���CYX�j�z����j5s��R��`쁃�i"hsS� n�sz���'��LlD���a�y�幁�����D�$�(J�+�F��k�#���G���	���2&���W#��ӕϧ'5U@_�TMP�n��》\����J��r:)� (_�5��ș���F#�<]�����Orl�1*#!����9=� 1ɦ���O8�f��ʥ�UZ�TK�������*$�CA� ��"�>��J0�	����PХz͛6l���l�.q�PD�K�b�
~G2\�D��˺�A'-�sv�*h ���掶�P��V�օ�\�*Te*㇪�P��2�A��L�)�)��Z*<����#��
�\�As�_�ߟ^�J���d �)�Eҿ8��0f���kUP'�,��텳�5�M�ct�@�<�UYD��P�ʟ�*y�QZ�*#��hGdR9���2Д⦃ȕ4 �S0�B�JySȎ%\0���F^�#�.x3�w�O�}�����(ʃamH�ca0���:,N��z��z�K%0���V6��7G������*{>.�Z��$|H�(_�[#��F��0�����"���$"I�CQ��w5�����H��5�%��vr0S�N".�G~n�s-$R��C��;	���O!����;��[�j���)��ebz��BH)+6���kDI���P��n�L�7p7�#�]��6����i��կ�7����$�����i�:��
#������ҦM�m�5�MMdN�J�$W�;�L�y!�|�X��-i\�xĚ+,V%!&����::
f���WHFԄ�D�X�I���7l�8@��!X�D�4��^����izB<��LmT���S+�MA%`չp����K"YzB:�'pjժH�<9����m�=9����b�oc =� �(b9����a��)���B���Dd��.��eR���T�ʤG qr�s(�@�U��K��
v{8��Dd�Tr�<0�As�Ueq�H"e�6hOJ$����z�cdtxljR'/���'6[�
��xa��iP�a��>0j� ���6Q.AL�e��R������hh�f�Р���<�N�q��R)�9�ٳ\��H��=�2r���%hAR%Ǖ*JЈ��B�]DeRPE�4�=�\��ѩ婒�R��2;auUY���e���i`\�Z34ǩBy!��?5\����E�tHLkL3U>�p�e�HR5���K�p�ȴ�tz��5!Q��mnJd�Z��H�>Y�T�@��˒�h�&,D���R��Pe=s@�aP�s��L����C"g�V/#���9�y����}"l�#O�7ɋd� ���`����x��D��`Gf�ɪ&ލ�,Q��ܣ6��S���*��PGD�x�S�9b�5	lZh�'@D��c���Ci_E0��  [d1pNOm֫e9���� ��a��9����Ͱ�1���6�e@����Ev���A�t�EJ(����V*�<�䨐hb#�
{Gl&(%z�B�C�CB�[,B�R$K�\����"\�A�Vl�T��J�Q��;BT�	R� ���&�a�n�vi�>���Z`�-�B�P���D��RV�Ǖ1rl�\����R�=fʂr��ctP��vW*D䞶nT`~n|���+E���c�z�As�Txa�*��Dd�Ah��g�-*�ct��I\�ҹ��a�C *͐No��.a��]��]TЂSȆ<0��Zh8e��ʦ�*��TЁī��Td⣉W8�bP���\�C�/`�#� c�t�1rh"}Nl	����M{����p�Hخ;��)&�$�S�}-~�#ROl,Z��i�jn$w> m@�9�Oz�	�(/�ѧti��ڛ�'Q�YY�W�g|LVN��.�R�������hV$��g�ZW#I��zh��o�N�#Q�����+2q��Bn^)����Mq8F�����:6G�Q��5dNH��m��� ��8�bS5���eNj��@�'$�ErE�4�I�*y�#�'3u�a"k����~?t5�rD�Yl��Q�Ė�&9:��"'A4�47p\����ݲ$֥N{>:�qr�?"t;6GC'.~i��G���E!M�j'�T�#�Rɵ���8��'>�	�W�zBi
�"&�M$M6��-�4�@�kQx��p݀9�(���~.����n�''��{�(��s��%2(�Q��hJ0�QG�8��B	Q..��hhG2p29��茞�B�.8yV�IZ<��*�1�!�eq�C��6[O'yi�I�R�jg��$����48��4H�HtM=^N�����?n�=�b�,���Cf���0���o��	R�6P�ٲ��r8aV[֛�$�o�Ӣ��(F��>��.�9��Pj�-�Zmٲ��H�Q2���.J(�B:Y�*�(02Z\��̹7S��GD(�R���2��2�e ���F�_}hl�J���S�F#Y	bLmI��ȤbkI�!֨�����p���m�|KI#��M�k�zF��#i�č5���3�kn�i��BԢb�#��sك�$�6~*� ��JB2����p[״r%;��Y:6���N/}hvl�&"s��I4:ߛ��a������dn��-l���Ǐ�4�K�\��y����U"�ʌK�i�՘�߷�ճ&Z��d��T̭��N)���"7 X����ș�aA��bqw�닮\]s���P'�E�ri��}~�A**�8!B�_��8y-��4(�Q2���.<�B��R��x�UIZT���6hh�d�s���Ҝ<�R#�R�~G���&Y��R&!Tиᔨ� x��w��F#؆��J���
}l�\���((  � @�9�����"h\�rl�A*D��%D������ےq�K�2d���ZT�RV�@�Ӝ�9�� �0�;�a����+E��0CT(��@NG���Lrq�q���㇬�0�eGWl�bHQ!hT�Ȫ�W*cA�MU%x�:S"�J���C�.e������?
2�ء��?
2 0���
G8)��L\yQ��OϮ�܌�O��l��7ĉ"�ȜD�4���r"i���Q����``�j�z�T�j�5�v-M
n�5VF"���<ڶ����KH)Ɏ�A9D�%�������oB�5�Y��+6�e��$�y�&��؛^�Tޔ8JA�H�&��My���5O#M	�D��jNq:/&���:���ZWRR$��h�z(R����$VR�$��m�8��B4�+ƴ.�Lk�ci�%�M�H�"n�@�:����M�����^Z@t.�&0x��Y#Iԅf��iO(Y8&���NNi��.bE$RZ�i�˴�:ަ��&�IbSRG��f�B�8����d�|@�Su�6ޝ	�y���6�"km�+M�D��A�����+,ǚ�zHҦ_��v��&<d�$��?#��~]�bT@[r�Q�U�P&`	�28�.n@� G.�d�:S"�#��PǴs��PJ�q�Ȓ�*2���9��uFR�"����"h\��1r�*h<�L\��
%�1�&2��4�ˡN�l��]���M{z�S���Y@�IZ(�0�T��lH��xl�xm=���p��6l�D�!��c����86<<b+�K�������"Av��Lٲ�yR�ʘ�������I0�&@���D@6�07On�S�-1@�PЙG.����t�_��**�.��98� Fh���F%�UB��b��c#WX���Q~E� �a���ڜ1+U8��y=�����L�=H���;����u⦛��z���T��9�_�Hܭ�V�=<�(�#d �`!�ad���s�����h�#�@Zb�������"Uj��M�6&�~��:��Z
�����@� �Ȑֲ��W����8f"�M�Mr����c9�Gr.=f�F�d�Y�7�h��0~��Lϑ��b���F�@	���q ���P��x�J����M�� {.Ў�B���e�C-G*�By*QG��9�a�*�Z+A��6PT����M�٢b&��L�f�,�Jp�q�lٲ����؆͔K���(�!ga�K�<\er�4J3�$ttw'!�nk�@ɒ��{{Dq-�6X��lٲ�\�Q�N!�e����ONCh<�B�2͚(��9��{rv7*}NrcB��0@����"G{0`I�G�@�QNO�3�45H��.ASB�0ᖄK�2�R��V�T��q*�W4D���Z�u)�E̴#�J0���#�J��'�Nn�� `'�B��
G8)��H���rPM��yЍ~֨8��5�i�eӇJF#��SL����МHZ�'=[Saj���+(��d�5�<�4vR�$��h^�i]�kT��D�ېͦ�h5�?�!��{(oSǍDi���5�O#6�����D&���X�����JF���cq�AXbKl��F��hj�?mZ�@��5l�Efܑ�'�)
Mi=|��Di��)�#�BL��y^�s@�j*tZ�SPf蓙��]��k��m�2�ڐ�v?::
���O'yd��')@�R���kLw�O��6���'��n��lu��4�	�P3Q<��RoHI��ͲD�[7_�)�ǎ�k�u3��)�'bE�0uHo���H�)���կ!+��5��^h$oB�mh4m�&	7��3x`6�hG(0d�'7g�N@6T9� \��6�y�@��璮vs{�p��"�\3��'��`�Ea�J��S��?>����Te+!D�4Lb�,�
����"\�%�1
��R$2͔M�T����R�(Xи��8� �e�~pP�/�� ?W 0� �4�t)��S�ٳf͕� ����1� �\��Е*�Ǟ�_KJ
�GZ�V��r�ħ�hm�!ٲpa�&YG{THFTHF�|�O?l�rs�Dxav�AQ�i�㇨���(�r5T.�B�
:���N$�D]�d�C��.A��t���'���C@����׳�a���
r CŴ���V��$G�pFE#M����	�dM�#����ka��Iz���'��l�<y�~�C��e)�Do���7R�s8|�"OS���B#�g� H��t���"��m�I~<�c)A��6��&>܎-O8|���"><vR/��� ԉQ���OJכ�T����2���G��.�F���`��ͦ�
����<�����'RS9��b{��E�w��R��`�N1�{Eh=8e������!]��6��E��2��TZ-v���~)P�M�ٳf�ٳeL �SB�6W*D�&Y�y+E�,B�R%ʑ ��l�8f�-�4	��`_[%��v��0F�m y-Lh=e�T��K�*\yR�ʗT��K�D�K�D�K�D�K�D�xat�L�a��@ݏ/\���酦��-�Zs�m���6R�� �Ϫ`�ܪ�Dd�p�����\�)O.E\�ЊЊЊ�S4 d�#�%<�)�G��Dy��*8�)�H��1���'��#�Jd��J�����;�u� G�G1�
���L*"N?(D1ب�H֍[��&��~Y2��o�I���NYnF�D�#^wS��O#J�lڦYǛU�U�B>y�ԇb��\��"m[sr�4�֎�H6mY�� wA5|bnHdI���|y��T�@�%�[�sx�+)I�g�����χT�@e���#�L[���v:�k�r�5)��F���9̩�5۠ec�A8x�[6����S�j�p�HM✤�;�6��bnS ����t���P�oI�%9e�O(Y	7�&�j�RVԵ4NR�F�L�S��$g@�zh$mT�e7����}F��œbh.�)�59Y�z��v���#pI��zh��(I6�复�L��;��P���hy��T�i�B�&?5�%rh��kB��r��:�&����]ԜD���BI$�X��J��?�9�ߑ�%JqR���T)���'�b��[l9;'>�����\ �!�� 0c�;A��G)��28aIK�AR+("b��& ���b��.A�hlB�,B�& ��"cA��K�Dк�
�=�Oi�9'��6[� yU��� ����s�2A���:=D����f͞�*_�  0`�"D���c����"D	m��_\��	�cd��Bo�` ��`M6�`ᔴ6k�8(a�A�h�֐<���F��?Q 0 d4'6ʈ�,�h]f��*�n�����sUc�uJ�T���!J�\�0a8˳��*-vz��]�M�Z�r-T�s��O�HƩ�"�{O~���<�]���}�T���njR(n���܏���c|PvkSɯU���u���'q���Bs�� ul���ݘ1�u��{Zl4���'�-�S�!Df&��8�˘����^�fR�=��)ڬl�Gw�6Ida'���!����\���?Pj�r/]��Љ��М���n�� 
s�	��.� ��/OhvI�N�i"�l�*z=�\̴-�\�\�L��M0���6 �01����ypGU<�q���"\]r��g���De#(�E�H��������dᔨ"e�("e�("b�H��b%�1�(� �&Y�eLTй)�ǒ�*h\��q�K�Jdʣ�Q*h8�(���h"<������� {\��Q��H1�s1�s"h\��r&�Ț ��"b��& ��"b�D�FN
�e�Q����GD��U�(%<m�������'�/�`�
��㇫�J�\�aVWT\Pĥ�Y�d���q�Z.E\�ЊЊyu*�<��U�?
2�(ɒ�%D�Z�TЁ���#��\3�qH��Ty�q�@��	�S0أ' �(�{u1�A0�L�HړH's��"��B �z�6��Ƨ��ރD�E2�����,�T��5�y�)�gt��5VIĆ"4��u4ܷ@Ɂ�ч�E�6���L-p�bE2ԑ=��R�1t61ؓ{T��tT��MJ�#oI6��$w�����rLz�-�58d�����ٴ��Kt��Ӡ�xړ���JD��!�c򐄐yVӳ��bL�II (�Y5�F�Q�t	)�ii�$�~�s(o��CQ��.P�&�����h�L6bS;ƭ����I��!����nKVAp3J��Ko�%^h^5���#|BPo��ͤm�H��B>)��-�^KH�[�ۀ��0_�JK�S��t!�� m���V%e(��F�!,JG�E���ȵ�b4(��'�j��4S!���]�o����� ��#�JqR��%\�(��'��`���2(�Q��h\eR#��\�ʤ��0P���?=�2�]q�TLAD�1L\� ��1rCCb!b1LAT�RV�IZT�q�GG(c�8g`MR�����Y�B�`@ʌ����A��.0͖! ��g�

s���i4��'��I��X��M���e�
��%ʑ=�~"(*(*<����aG�PNo���49d���bw&��$��gg��Ϯ����n�80˲ۚ&��*D�+B�PУ� 0#i��cE*�<���ǥ� ))��.�i��#i�Mʊ1@Z�cԡ8m��R>A��(y�\l�����~F��B�\P��!!4r�hH�jl��� �<�nBXϚMk�&Cu�G$d'���QޛX4^'eɇ���D�w%Ȝ��h�k�N�!4͠v�=�,����tU��˝V�h�PG\М�~�mI�ˡ0P���M+�4���j{)�R&'5�M�&uZ��� �yl�m�0��M0��?!8�v�(*�F���[U�s�t�����%P(��0��ؑ�e�D��-8�sA<P#u�B�6��BT!\��Y�V�U\]r�맴U��*��EhGhT1ULTй��ʑY��*�.T�LD��Z*b(� �6l����!f͛("b%�1�-�#��r�G�8pP'�KnK�%�\��R�4[r��ɐ�oc
�B�
�+��B�
�+�����b!b�'7�g�!���~8�*�,�4%�e<����m0���H:1�کr�u�������&Yb�Uer�G�<��͓�ZJ�R%K��W"�E<��S�D]*�H���\b9���\�����"2qR8į�
2�1)����D��!H� q*��>�~�q0��@�z�G��d�GCt��|:�LY4ȓF�Gq��DH�&-���LG�m��Ĝ�l��u�~�''���ϖI�f�Ց�b5V�V�#aѹoT�Jp�����mMm�X�RY�K]�׫ZWRT�������q��p��f�!�R��m$�n�h�O�F��03i��`$wyW���!/��2�L�:\#U���F�[p3��iY�-Y;#M���Y�l�@w5��K�1�l���m�ĕ�=8��R)��ԃV�����5 ��A�f�IV���254W(R�$�S�Ұ,��rZE�jS&���6�~t47D�nD�r� HĦF	� �h.�:�eNf���d��2��Z�E�zE��� n�:"}@D�L�q�b��9�0m�{?>o�顩�#�Qw�.J0�ǱG�
G8p�A䫎h�\�gg7�7 G��%x�:S��O#�<���a�E�����������b�%8ySB�1LAD��1r\� �44L�e+�b��&.T��T�B�"AR#���S��F����4�O�M�3D�6F?#��1Ѵj��� ��f�CCGvvvt:�C���� !A�'�	��в5)�	�.�D��6O%hv[s.(e
R���٪E<�+��r2�'�$ެ��B�##Ol6�8&:D�-7J\�W!]��@܀��b�Gl>��]��hr��e�R�hEhD]� ��07$uh�Xe��JrCu:5��"[y?S�`�̖�7�Vü����	��	���I�bS���)h��b��L�XZ����Q��~Q#;��lk�7OӔ�Q���G�ʭ7�M�"4�w?;�&ﵳ�n�ku�_���s�u�L�`ƛ�d��f�M���\���N�@3ef�x����"��M,U�ȩv�������)@f9�D��K����sF�^��ndGw{��u$���Ug��&(s}$l�����&��V�����x���s��f��E��'�<(�#(��@�#G}Gb����"b��&Y�e��<1����"b��ǒ�.T��X�SB�!�e�D�6PD�6lٲ�&"\��ˎ8dɑ��?  ��,hTƅE�?�涶����*W���  P�������ٳf͛6l��q�S@�댜a�$*�.\S���A��H�ޕ	#H�F	C?#��<0�&��L�AR$K���*�.T�͕ʑ*h\�(�Q.���R�Ƅ�D]*�LJy�-K�J0��t���{G2\�8į�0 a���J0���Z.�B)�aA�bTHS��HȐ<�q��Nm5��NI���%<�B��:�%���m�k^�`�l#N�N�IRH�}"\��Tt~7o��,[�R[���&��0S��A��wqA����"ڈ��pjL��N#pԅ���Ę�,�����4Nj�5�r#}l�P8)��n6FH�G�dP)�	]��mѷf���~VoIih]&�18�ͭ�h��6� gu+e�S5�k�ZWI��iִ�H֛����Y��1)\����Z�p敁����8H��	�u�Ė�&���9I�)���v��H֛�4�1�U~N0t�5�Zn����������S�' l<��)ӈD�Yd��w����&��@ڧ$�6D�?�|�<e���t�%utm4n�;���A���J�	#K|Y4)͡t��
q<T�͒2��@'&�r�ܟC8�bQ������'�b� G<]�(��ߌ�{GG(c�9���?80�qC�
�0�(�Ҝ<�yS��
&Q2��L���e(�\�D�0�V�6hlІ �����ZF&|T`�>L�
�*��Y���y�$ښ������ݞ���<<<׵�z�zb$LD�����M�^w5'�[*��\q-�FRٳd��.j	�͖�7�q2�4.��"8ɲ��z�F�!��J�.hh����$z�5KM�l�.��ꨫf�E��ȵ�y�Rg��)�p���T0�B9��(^�+`mz�3U>r0�l�d$��*� e���-�U���쁫OGR�/R������ԑ%���ף\��ʛ�⥂iJԒk����)��%f��hl�I1���`mFώ[	h�.e�ڱ4�+���m��٢���6n<56�0P[#>[l�L�8b;e�����*/(K"<0��n��kZqԷ����=U�V����h��@"�.��O��8`��k�G��VŠm����%H�@Vp9�&L�[� ��������=�+�Ug��R�s46l�8��Y]��+
<�b���=�)�D�7#7 �quˌ�D�1���r�R����<{�˗"D�D�A�K�"�f��\��\a�ʑYb�2��,�<x�r�D�U���F��涶d`����@ T�P���f͛6lٳf͔44;=Sʌ��B�8'�����g�(�%�<�*-~rsD\����zrWሒ�Y��R%ʑ.A��b���;,B�&YA��Ub�%�ʘy��W8��Lh<��Uʎ.h2��:R��L�<�1+�!���~.�(�8ģ��\��H2�bS�W.E�e�A��	m�S�Q��mbp�W�֙���?6���T��y���V7w��"F���M�<V[F��ȍMWy1�47F��V���E򓡭5��Kʔ�Ou���3���!�~t!4�����͒�bg�{ս����ؕA�8��<��@>��E'��9�e�+���ӊ�mkr��΃H�����Mbn�#o�F�B�NKH�
�'��J�+8��E$ǩL��K?yԅ'Q�f�kM�k��KH�Ii�h$�j�	�
AZhu��%sU�Lv(kѫ"{^R^,F� 3knW_Һ0xԥ*X�K^D���JySz��_�7R5T�"��5HRuI�ב9̵H��S���u3`�Hn$��9K��KE�j_��v�^�F��F�N* o��T�u2�Ib5oM'b�	Ĥ6���=�.e�*T�<)���%��g7�b��J���Q4Tq(��ˀd1s��O#�D��Q��2�\��'��\yR
�1������e(�\�D�1��6lٲ1������&_�̿#�١AR*&.<���iQ�4�u��PD�����ڭS##�?;99uFNW"~}���vONl�O��*�W1qt��Dd�B9�I�ED�o%��dm:96T(hL�#�ۤd��0N�ʏD�W��R'4�&��:'�Zlh\��ʟ�WL��l�6\���L���𣊋�48e��P��#�j��D�ک�#-7����� �b�r�](�}��UH6��n�s2\�=��Dp��P�l�5[��r���5!55������*e ��$��MU��a$~���A�#j��R'i��d�>�^Z�$}vh���Lv@Uh�'{-O{PA8�V��˜�L�< Sz�2״˖O�GپHx�zٖ��L�`��mx��b�JD�(G��� D��'#-�B`IN�)8-��>~<~+LP��M	�ZEvOR5S�Gǚ� �Z\R�,�+�T��U
;��W\ĬT1Q�UU]��W\�0l�K[����8�r�H ���b�˚   ����c�*T��U4.Tк͛(� �&%8y�l�<��)��"e�6�˘�tH�*<x`�I��ttqB�"D�����c�"8�R�͛6lٳf͛(hhhvz��cB�FN6��ݔ�8��l�\0�r+$BC�������Tr�l���B�p�B&Q2��L�����1U���1��#�W8��U�̴2�y*�ʙ]b��L8�q����h.e�����Z�Tq*�q�^�#�2й�2!3ʑY@�T��nm���Ct�ޠn$&�mF�CQ�!-�Fޞv#<�F��p5�kp"��`x��)�^���"i�ȄD��LR#T�!7�0�+���ah�X�����d�aRH��ڽ�F�O��Ѵ��t�qTH�`��=F���f
v��z)lMp��qȩ�j#X�S�W2��u�4Vd1��"�m\K�ԑ4ll���ed�ּ��NVH�
JƴD�6������\4����T��\��D�k����)��*A����	��^Op�ƭ#�ґ��%'�׈��!���'��M��H.�:w}6����кL�lF�����fn�'I6�8T��� 5<M�? 1,��'b�>�<�e<�]A�ڔ��
B��^�#ysL�ZM6�n�P�Z�ctLmbׅ��B�$�4@�^ˣ�8e��0�7 Ki���oo��.x�U�ҙp`b��{G��1�c�; ySA��4<�+B&��\�����
&Q2���1LA,�A.B͛*��"J�f��S��"��e�6Q4.AR$0ᔩN��3�%J����%J����Щ�
�Ъ���=@��ܨm�G2)��S��P�����j׻�.��Ӂ��xa���P��)X����.\�6R�8֚��yݵrl�1**T-����_�N �3Bኒ�%hz���%.p��,2z�]�Pz�';�.G9%<�^+}\)�8D�l�"Pk���4�j�0[TP����)b&�6�".i*kB$�կ)����a-ش���l|Ô�rbk�$�sJ��<�V�nv��v�%Kb�Ei"(/�h?r8n��~�h�ll5H��6ü�r&��v�rS�$�t�@ڱx�[�g�b�o\�ԩ&ɱ7B�~�#��*{ :�� n�&�O�Q�I&������7[4��Ĝ۝ԭ�1UAsZ�)7$�SM�T��g��boU���D�X�5��kg��r8�u+-�"�T���#Q̽�T���R��$u��7f�$wb�Z�u�R��ʪ��C*h\�/� �$H�8q���+&K�{ b9uʑ.T���M�ٳf����rS�� ��?#�����^�5!TйbS���ҢAV�f͛6P��2��L�eS*�T�&Q���448p�:8�����v���'��MR����h1Qs&C?'7[(��̿#�9fɒ�*D���R���L�.D�R&!b&ZheV���*#�W%8������.y)�K�1�X�S'8���FN*2qQ����Td⡅�2О��Z`~��M���t=Q�G{��ur�N͗�j��w�	�v���:��K���=��[����hDD���)��РHY�p9���R��S,MBD��!��t��|�2�:]����ENm2��yHMz��r%9-�6Y#Y�ƣgE+jO|��BH�':��F��AĲ:�1;͢&�$����^�h]�Z��Jj� H��z��W���;���E���a�4KZ�V�59M`6��Ԅ'�u9t���ZhI\Mi]&|�&���j�NRin�|o�K�I|�1$W�&��dl>yČM�5XHViA'�zܾ �j"6��@YR�Vo"j�$KmǛR��м'8�i��N5i ����wR����Bkrؚ�I�6�NŠr�nf�䎃�jng��ŽkJNi�bF�%Pr?I���G�����qF^�?}8��⟋� �)� �p.d1r�#��S1�r�"JЉ+B�"h\��Vlٳf͛(hh�D�&W ��1r��&.T��lٳeʨ�e��؁�ښK&��Y1�f͓�R���Z*D�"D�R���3�T�`�M	R٪\�e�%�i�O�������MP� �o��J�#�~��5�o$ґ�AmPÌh\��L�t����\�SB�M�֛�b�k����s���E�z��{]��x�:V�ȅ?#�����9��{E؀�~B5 �=T�zg |�D�L~7m]���(#�V$�M����Uͭ.�>T�Nv�Z�hI�koV�2��u�[�z�o�ܥ-r[kޥ�&��GF����d������)�D��*LoD�l
D�2����n�hl��'��ak|<iqm0�>}\|�n��_���kV�I&jK-<Yn�?�/W����Iw��L�&��א"憙���L3�A@�D�SG4�9��Bn�i��p�<��6�|`�kׁrs�ض�j�"N:$DC�s��Lt?mGC9;��n�A���d��� �4/G=~.]����r�ˢa�Oh[Ls-0( -?"L8 ��]��if^ҽ�=�<�r��c� ��"A�1��$H ����M���z��`��e)�VU4 ���ʙe�� ���ce�6� $F��[�0a�*<���U4.ChA��ٕK��*C�f��L�e(�D�"e�19AA��4�3�ۓ�7eFNYJ�0���#?(0�]Cf�e)s�i�Cˡ�D��H�2�4T�yR��,U�2���CA��$�2Д�#�W2�d⦃ȕ4 �yS���%G�bTq�Q�%GG<��x�9��VZm���Ԡ�O���e�
�S�̀}GsO-y9&#@'����54�:;5RKbk$jȤ@ޅ�^Eb� �1~M,���&�N��%8]��&��%cz5o�P͇�#-U��C q�]초y�hGL �G2�(z����f:�&8
i#Sn�)8S�!��fF�n]���dF��Ԛ�mM����&,Ԅ�ݺm*IF�ʴ����ccV���mm�]"% I�jm�"F���<M�L,�)�I�f���@�
qF
qּ���GBz���|,JM ٨�iY����"b@��%5�'[d�y��{*m\��f�ԥ�M-�۠D~ީ��%q�f�y��D¥��NK$kB�"�n��C8}#:��j���S<�+��Ŀ,�����d��6�������z5S�DKi1(+�bbOn�b�I_Kg������ѫ`��� ��+A���Gd�Ĩ⌾� [l9%yq�ˏ*�ET���Tqq��� yR����*JЩ+B�ʗUf͛6lٲ����L�er\� �!TйL�d�V����l�"G{�`��RJE9,�NY7��{M@P�No�Y�Dи�r�l�JyQ��K��<0�r+4HZY�D���t)��I��&6
�� 
`Ô����ZiᜟD��m4�w����6�������p��۽$�0"(z��Ĉ�@%�˪��2��OQDd1s��(U%hsNrTe-s-�UY�&�ې�V^�l���t���"� <��ψ�k'%!U�� 57��2���$:	d<�&��#h��T�$B��!�������D�$aPnbY'5�&�4� L�9oG�ޢed�r�jkAO"�ٔ�:4���
 /�`�P�������v�^~qByq���a�00Ե�Wr'�7Mn�p;7Òxb�At�t���M4�2���x�R�	�<$� �Z�h.vsX)ӄO)#�yM��NI5	�R7^�M�E�-QNM�5�ޣE��l�\�y*�A�=�1��W#��.PG���\�n���*�k��Gv�|�ZHTPF�~�.�Ͳ�� ��p������@��ʕ*T�R�Ǐ"D��1�c?��("пH@D��	�8�H�7-LTЁ��? 	ءA��2Щ�ʑ ���O[Nr�]Lb�ʬٲ������&1�6l����Ç.]�S%� �SBsM�h8�c���$��ge�'������(2�ЈS�g&�s�p)��ցG��UL�"CB�>�(� �C(�(�Q*�UAuԩP)( H�!1�$q�"����d���h@��B�%�0�p���x��Cۘe���s���C;9���������nD6��"L-l�����GA�E8�4�6Y1�-h�|�m[ƧA5�BuGgX�jnQ�kxڕ�i�rD�~Yj�5�Ș]�hr\]=qŻ.8���#@�yw�
T��5��կ�:
b�IčkU�Ks*oN-�i��M��j6�)7�ri���x7�uj����mK�\	æ�Eyh�<ڬ��yj��w�S��Ū@h^k$Yѩ�����I��!���\C����bY����zW��c|OI�N�kr�_��DJ@����DtS;ɪ��KH&ڸ��eA����&1��s4�6�fԮ�),��m���bnZ�A�),Jm�ML�S�[s���wY����F�c���T�F�M5D���O�n��۳L��Ȣym����}?��� �z��,��	����R�h2(�`����Е�W%y�2QH�%�]D�*bSȃ G8��)�Gҙ.q�,�b!c�1�c�1�c,ٳe�X��PD�!b!b!b!����Ǖ%.q�m��=l��z٨�b,�J��1b޷ ��\�a��젞��i�����#�F=��BЩ�R=�U��Vl��U��롯oIerzh�jn��99�d�T�0�l����	��S���5ȭ
��a��N?;>�#@Ě�dC�P1�x�;��s
9΅���D��E�
2��\�s'�Z�Z<Hד�*CI��H����(OoD�	ɢ���	6�6�l�۷I��d�tX[&�;��M��_�X�W	
oQ��%$���hJ6����m-<��jb#w;U��N:�6�һ�-W�DI��\��!#G5�뛼v�[Fnt�ÚV��_� �}T��$J@��"�*�E]r+���sISCj|�"N��!��zPBy6�k�CZ��
DP)�~�0/_�n���D2��ӏ>���Jw��Z@x�&�R(=S��Q��%8�5N�F�~�Pv0}r*s\��{�su������P��M��Q=�� 8�����P?7j��l�̠������s������q�J�*<x�&Z?c�1�g��6hZ���r<q�7##��HuA����J��Y<���0�qC*Ef͛6lٳf͖!�f͛>�t.Ty*�1SE�W*~}v ��s?0j��"DxP��*�G�aÁ��Ov[LN�uV�.�E8����˗.8Д��X��LDy�P��X��T��%J���J���
�0c%˪<y�˪rr �n�''GG<q�'�8��`	E J���H��8��PNn�@-�94Ϝ�댿4ό,hh	�@�@���@uqvȧ4k���\���l�H��5&tL_�]�7��Dכ�d�c��]1~�ww�B��	��S�yB\��dD���l�3D�<��X��~�F�Ƥ�BYS��T�)�W�5�8�~S-z���D�#��^|Hڼ�&��I�����]Ԙ�4�����f&���6�Mש��bLp�-�5XT�����m�<��L(t��E&�ȜDwY���=x|ބ�MGb6���4�ަ����$VX)	�4�	�Hש�ޤ֘5�Si
��iie9�Z�8V�&�$��'��E�rqS���1�E'��zyzZ�1/��A���:��ʙ�i5��B�#J��H�6ֻ�R���4�V-2'A�#|Z@tF�MI�I$����Bh���&��V%bF���,��7Hӈ��;4��8)���'��D��6h��� ��1�R%J�4.<Ё�"�A�B��� �d��K�b!b1�c?�͛6X��X�Lb!b!b!b!���Q1H��
G))s�� ��|T`�5�Ci��nFPЎe�
�8 0e� J	�����-�7L��}l( ͖J�)�-�7G������;��	���H�})��'3�%��PT$�p6KL�-1��٦��
͛5K�('�����A��I�6�_�N[�DÉF=�@򣂆49CDÂ���B9� 4#��\� ���˳eA�����C�S@g�k!��m3��EJ"rH
�I�ۥ&����Lo��(L��ht�D�nv�:RF����i�Z�������7\�m��A�G_�*l����&"P} j���%�x��gy��� ������M7k�V7^��
���;����F�`�U���SU�7R'�)���ג��@kkڣP1�����v�k��0��z|�⢑� D�d.;G>+$�;ڱ0#e��S�����L��Mp�yr�Q�1�NN�͔�3�H�%��5C
 n�i� l�R���[B��6�y���~r	A�m19m18��z+ �����F>��9Gv�1��U"h\�R��0�È �c�1�g��6PETЀ`��Yh<��Q��MSt�g7��WY�f͖!D�2͛6lٳf͛6lٲ�,Cg�J�'(((7S=�.���'%�5��4x����(#�/��=A��Nj	��Nm�$��{�a�`!K�*D]u�U��hhhc�� �s1�D��Q4\��$It*�ND\��&W%J�T�8���Qr�"�.���@llL����Pa��#��e� �׳ �#�<pR���0���9�6���4����ͺ���\0�q����G�-Q'f�7���O*R/�i�Mk���4v?p��LI�RhY"`�@E��@��6H 4���Nj�V-�I@��<��D��<�;U<�H�5����m����Q590�bRMv�HVH�N��ԑd"z��¥�9��4��$���bk$���|L�A�P�կ),���^"H�	5�����hV�����j�o��s�ĥ��$1�AG'���9"Dt	/Ʃ��Z�y��K���H׷)��su�N4�SGg���%��K�H6VZ��[ŉ	�$j6&6����L5��i]NY5��$�^KH�7���F��kn�0_�ϗ��DI�4ЈMbNpN�����C���֬[Pi=f�46���'��bjw#�j�Ԝ:�(R���i��5�1&$����
~\yU����U�Y�\�Sǎ8e)����Ty�W*aq�Q�8e�SB�ʑ1����f͛,B�,B�&1����\�	�)U%h�DƂ��^ʇH��'B4H��t�t�m~m�ɺ�#y7�&����u�:�n�������Ze�=��\���O���!�ѽM6�ִ�Y��Myd�<�_�/���4.�S�E#����ִ�i1:JE#^tw��I�� ���SӜ�
�E��:Hm��t<���&�aĨ�%8�*��)Q%h�eQ���Dd�#'�;=�[vhG3hEJ��Us��&y%z�g��|��r�SJ;H�SV���iL��I
#@t��ȩ�it>���$��;��DE����m�ݡ���<|~tvp	�n�n�&�q�2:��cu�N\�[O_�?�0hLOT|�:n0��(l�b5� ���a�Qka�A̦:nWI;FߌDke'�V��SZT�1-����i�����r�'���#$	葮q��3Y��lp'�E#��j�����{z|�m���Xmr5�*�rgi�}y5V��IJ������&�y���֏7Ji!�{jFRoZ��������~<��qv��G�.y�-V���ȋ�DeR"�T���FU.2����"J�(��8�3�1�c�����ʘ������'�Y��S%\�y%�6PD�6lٳf͛6lٳf͛,B�r� �?��L�.1����i��	�#IFď�H6���&����'�5��T��~�i�6V�)��.2��*��hGh��0`Çl2p�Å�<��r��ʎ.Tq�Q*�J��+��\�*�1*TD0cB:9�ts�������-���0	�͇0��M��I�b��{{� �g��[��	���-yY�;���#�9�&=Q[̹����)��E�^t5��741���e��y��`a2��ֵ���)	��\��L��b�ަ���C��b�#Lu�y5��q#��U�H�)[s7S�Z�ah��6q8���RF��M�i��@bj�F��f��4�� 1'��H�!u���&�' j��-�_LF�m�����m� o���j�T�@�~�I&$��Eb���:�'6�s�1�|Ru�jשY`Tt���i��$Sm��n!����&�BHӺ����;�I�f� 2i�$�R��䀦�/�J�1�H�%���Bh$�tZ��'#T�'�Ǒk��`$w[0S��;�O��o"��f�;��k"b��iY��N��F���Glh�G�6K^K��5�mI�nH������Y`�"YD�Au!L�t)��&'#�#/�g��A�(�Z-	P��D��ʌ�8�(� �@#��;
~.��K�"�bM�D�1�c���f͖!b!A��X��X��X��PDƃʘ�.A)s���Y�b�N�$0"(0"(j��;��ӹ��)������N�"�Nםf�3q���:H�w��JGz�z�T��{ԈHx���I�"�'Cȴt��`nT�l��[&�T�i�ri�,�"<�0�����M����B�H$�y<���d�o�K�zY&�W�;�N�t,��N��dݪq�R#�Z�ƅʌ�\p�As��
J�1��Csi��[v\�fyu�*���m����p�=����9RG�	�q9bZLoF�i�1��bZ5k��Sͫ��ji�bI >$|���S�������i��8���\̍�i��H��CmU ۰�dSU=+M��`�6Vߊ��]�j�6H���'��레 ��0H�4svĨ�;|~y�؎�.�L t-NmGV)��Ƞ3ղ�Z	����W��n��D��c��Xi p�Zk��tDN�F��tQ	~��k˩۵�8�05��q���L~w�N(*$ND<����L)7�f��u�@d��*�]r�ytU�5ڤU[44L�١�]�Dƅ݌b�˒�J����AA1�c��ٳd�V�2��� �&Y�eL\���˕"�f͔1Lb6lٳf͛6PD�K�b�(��"D�R��Z�\��w�����1�r��r��N͓������ۚ�{e11��i�6�9��.z��䨨Zұ�s9'''((9������ �ᔧ��4D�*�NT\��&W<�J��0�uO���T��1��� �%~~8 w��*�';7S�S��>����aFF.����g6��P��ɭt�ާG3����晐I���ˌ�4��K$ӱɵsLn�SO"ɬMdh~*6�D��=h�!?Ċ�� �������F�ŭ�ۖ���W�ԉN"k���؍dOn��7R@��ǩMNVZ�)�H�F�ڪA㡰��BI�����Y�j��7RG�Rkdx�:�'�Im#^W=M�ɺ��`�4�5�����:�GO"\ ��b:r`�����e���m+��ԛ|KH��$�YJw6:΄��H��:	m�ZvLS���SZ�.�X���A��S�ǉ��Oc� �Gu�ԒV��9�5n��F���+��yj���oM�#J��j���R�$ک�=�0a�|bSJI����akȜք�i�"��.�$�r}��8�����G�\�
l�7���k�Bn��S���s�Nq<�и�zN-kχW��ˣ��G.x�%J�"�]Au�1U��Dиᔡ����P[�i�=�~<�r%�6l����"D�1Lc��f͖!b!A��X��X��X��l�h\�&"\���OKD�"(#l��[����r�17zIК6��s�|�I8�
��d�P4����Qj4I�&PT�-#$z���ּ�N%���#�Ԧ�:7�C�g��?U.@�E�4��)��ۓ��$,�.l�:���$�I8�Cã�O%� �4Hy�S�JE:i�t)#oP6�T` �K��Q1RV��� ����������������;��oȌ�����m�!�I��j�O_�;)��Q�"k�l��I,��Ef��AA�<��_�*i� 7sI6BM6�������	5Q.D��:Ӧ?
 n�Hւ�$�	���A9�M�*[~�<�9�Q�s���rV�x�s(��m�M�"sj�DH~px����b�k�L5="'�ԑ��e��#2`쩺�vh��<~	`G����e�0H�kU@.@�&�`$ݦ��4���NE'y�4�a����Ƞ��$LoGS�增������z:�4��$����գS�m|62�&�%Ef�+����B�R$*h.pࡉQˮ8yH��tAr�� �� � � �c�1��L��&YD�2����r%�Y�f͖!b6lٳf͛6lٳf͖!AD�&Q2�z4%J	�m�A�dS�Q��i�	��j�&�����cUm��\p���������	��S�;B�YA�ʙB�aÂ�%G. '�77ggd���7���8y*愨4%AZ&�:9��\x�'"~~8��)��S��g��A�~~8��p`Ƅ��O�Tn���;�e�As�K�/b	���r!���7f�q�y���T�\ �+���{TxNwNn��Nn��2��D�&����5������Z�)���~�	?�D�e�|�)5RD$�y-rs��M�j�
JBb���&mi���$��`$wX	���mkr�56�Jp�#|h_��r5�5bbH���չ|�Bki��IR�	|ސ���β':�楚���$Y�[щ�Kg��-�h�?�\��0�Ht)$Jm���)$��ƨ���x��1,�o��MZ��T���H��nT�׊H��1$�'��j�*MʓF�����,���[R�b���5�}#o\ѭx�;�^~����hI&NY��JcϤJ���x]�t=�/���eM�jܣZ�BH��"o�BjA�ك��4Oi+"�I��mu��$�yBI�:�� hr"NF��K"[���@MN����V�K\�RV�%�?? �xS�@�u�%J0򣋚"2qS���'щ�a�2p�A䫎h8e�r�Y��yR��˕"D�A�g�lٲ�,B�("c�����!�e���IZ,�rhN
��O7*y,RGCQ�$�)��Ll�m��# *F��=@ʑ��Q2�O��'-��	�<���z4H���j���
�D�Q!f�FN	��sSe�}f�,�>*-_��N�"���t�C��{e�|e�Q��ܜ��m�d���Ϣ�=�3A�ȗT��uR$*Te)��w�װKnj�р�1*�%U<��hD��2y�[��\����6F.7 Dkd���ۼ���~���� �MQSM���~�y&�!�ר����m�{e��^�y�m�~�$~l�&_^��M�\Țo#K|��]r#-A�V�pb����7_kfg�	k&��b���$i��8�L�@ 
	KA0{.T�vhhPh����቏��	�	��L��BZ�h����ƣpI$�}<�@�zT��ŉ���0�r9��Ԩ�T4������ɔ�_�F��6�L(H��󀌡�:��-uq��3��r�{���L�%Jx��w�����og��.A� ��Ǐ � � �1�c��&y�Ǘ.\�1������1� ��͛6lٳf͛6lٳe���e�44b$Vl�SCA��Q�'�S�Ȝ�-������QStLL��}��?;99;;;=�(aq�NT�v��ur	E#�'�=�9�8q)�"�
<x��g�C�Jx�B	PJeq�꒙\p�"���\����#��  ���������@�#�?~~8 qB��<���i��N)�bT��<y)��_�Č	 ʞ���BI٪�GPF��\���^F�5���Z0�]�T�M��%�1�bX)JA��kyč*'�5D�kT���NKQ6�7y��&�'�[�;����a�L8��v$�	��թ�7�t��QѺ$S#X�I�@�|Wz����$ޕ�&�U�5w�[rA�:�WyY"�'+	n *H��o���x�*eh���Fֹ�
�F�.�T���#�����6ԉHL$oB�B��u(η�\Y���Mh]X�+⻭bhu����CZ5�H��M��5bV��n��h֩�N�H�'(��{�~SR�;�%�rZ�ҳLw�^��6�$<ڬ�Ee��İ>,��:�`j�J�=�?_���r���x���bn_�����|5S�䳡1Lڅ�u�d@�4��J�OV�0�4T�,�����p�z�;��Au�Y�[j������h \a�f��r�xg�ǀ=�G~8]�4� S@��L�\�Ty�F4G8��ʘ�S�<y+CA�J�"\���6lٳe�X��PD�!b!b!b!b("e�'��*h]f��ʕ%h.(`��ϯi�Th�B4���t�Jt�|�y:�7C��9m�=:�.���PLn�8���<�x���44tJ�
Q��1b�Y7��z涶])�?����((7O�����Ǉ�)��L�Ar��Ar�J�t.h8yB�.AH�<�V��� �栜��Z*��R�@�B���݆9�v7l
-l5T�	�����"2� n��[�����z��;�i�''�4h���M7$+h��^�;����z�I)v�l���g.m�"�����-W�j=q����D.�̍�)r�!��ձU�x%U%D&����\H؛�݌�n��݇Zkci��Q���WQ��"�v���1��eΜ� ��˖��r�ZDKp9�6L�G5!C�ɪTލ�W�K� )��˗?~2|��4̰�5�^���*].�c�#��ǵ�q@�=��1/�*T�ɖ"E��ǚ��*T��.AA�"D\�tH� � � �1�cΩR��1�gT�Wc�r�H��$H�*T�&.T���M�D�6lٳf͛6l��!f͛,D�ˉ Ěg�� Dy(7 7C���J��99<���lm�w����\|nn�j�_^�ߑ���%G8��愫�%\�)�Ȓ�. 1�Qi�i�;��g��O��.e��B
�x�"��ߎ#�T�p�!B��d0c!�{{;CD0c.��� .]Qr꟟�]�b� [`��q)�ǎJ�=0������#�rs>z�&���m���$A�%����RM�$�`�?'-���	״���Cdl�D�D�S|"I��+S���4O-I����.�z��mW�,��S?���V�����т�L&tX'���5�\a�h �ze����>)��SY��S4�Qd��$X��B#���j�����y<�d{7o[�r�$VQ)	��I��ޅ�*B��~SZ�7�v��jT��	��Ę�R����$K"o�G��K��h%a1����Y>l�>��5�� �Xio����[z���*&��Jl�A����S^�I���j��lҜ6wF���&�D� 6����BjE�Y8�t&��ֽ�n��m��\�n��t��G�Fבܮ�;� �-��	�
B����F����5f�oI��"�&����0�H�"t�,�	Bo#Ȧkw��p6ԮF�);�R��ٴmbLl��ɣQ���~��h2]0����Ake��b�P�� �Pc(����.���� �2���A�K�1SB	N*8e)�)O%hh<�r�H� �,Cf͛,B�,B�&1�������"\��p�V�ʬٳDĥ�%.qV��'f�T�m��`D&�y7�k^�p:M�ȴ��͚��l�!f�R�4����m��������R4j5���		Ʉ��c\���441/Ax���*T�R�A@��
~{�����`ゆ1*9{5�.��0j-��C��tce��M1�mX�L[2��Mq�Z���M�~��J��|6�������@#�5��.LPI�#}_��4��4̕-�n���sh<�TH�7~D`��T��1��c�tŶ9�}(j�l9.N��sK~���ǉ��{U)R��+���[#Ne�igl5[mյCL��BЄ�'�b�ӟ�����V�˽=���2�)*������)í03k��l3��%���K��5]�k�(
\�3KD��ry-R�%� �T�RT�R�J�*V1�c�1�c�1�c�Ac�1�b �%˗1�c�1�c�1�c�lٳf͛62�(2�(2�(2��,B�& ��"b��6lٳf͛6l�2���0׳/���*2q����T���Mm��.�djMS���Nnf䄃���ɾo�

Jx` ɇ��NNE�\���J�r���Z'���(6����m���ܜڦKno`�
\����<ÇЎ�y�CE*T�\0c@�IC21����4Q��  \P��˪GG<��1������uIU@����H� }k�#SP��JM�7�Ų��&�m4Rs*IL�r0I	�CHI~ޓI救YL56/���z�:tP;����[�"6���%���W��ud"_�ۗ�jloB@fӱО��)�D�'�"bp٤�bh?S�����`�pA5�"r�rxU�5%�хN��Dj&7��ZD��imՍ�
[�̍bM	:�k7��H����Q7 ]~wq$��m�]NR_<���u���U�Oz����LJ:��&�����Vmʛ�a���|RS?�y=0u�"I�@�2���n_��rjR���$���LVJpk�b|#N����"M���x-��xٻȬ�P�=�)���F�D��M~K ;����ke~b;����Z����#�2�v��l��7w��&/�E�����jU�y�b�����<���������5!�HBI�k"��M�Si�,������8������#�G��tO���=����K<�0�av%J��IQ��44Z(��?\�B�%<���E̴<й!��T�͔K�\��'��YD�M�*D�&Y��(h�AD�1Lb4,\��ʗT��r�ʚJ\�a��4lm~�t6S� Tx�����%KAA涶�t:�cm��e�~~T&&p�v��J����#�N�[OOhJ���c�1�c�1�c�1�c�1�c�1�c� ���g�'f�cd0 �* �����o�k�@��O��֭�*�UH��r2��Tޔ�IV�;�����Hj6to���I���ot8]'��64��S�;���ؘ���"\`��"LRS�1<cؚ��S\����We�R&�g!��#�r�"�:�1�M��=a���Vȧd�d�<�X�����ų#��7��C�Q�U���(&&
}~��c��[}}-n�7Q���5@=��
u k��ʘ�38��l����,�s����K�EE7^����h�OFZ�pP#%�*\��)��GG<��r$H�� ��.hhhhhhhhhc�1�c�1�c�1����AA�c�1�c�1�c�3f͛6lٳf͛6l��
��& ��"cٳf͛6l�80�R����	�=l3�#���J	m��A<3����>�M����-��|�5H��f	��nNh.\�1$K�A�T��0��g�
�
e��L�Ht6�'�
�F@6�7>2\񓊒�AR�CE*T�\d��8�ɕ�˪1��:9��T(RP����x��A�È�By, �l�.\�8���(5H�B�|i�s7�9���%��Щ8�&���BI&�-Q�5�ڬLGf���t�n�gC)���ȑ�f�+8�SD�%�I�Hm@C��v~Lw�&�<گ��AĜ�mJ�$���W/ɣ�+"�����1)$Bp��j!�Q��+�ѧ@�^Q��E98�t��y�,�H�i-�%���S���jpSȔ����"kT���"���Z�z�F�JR#i���m�E$�Y�jgu�p4�[�����@�i1�c���d�=X~�4��\�e��5O���l=T��Ș��	�����N�Rփ�t�j�;��;�j�5���\ce��F��N��5���$���n�ƣm���Գ_��ň5���M�A���	:�m���MbNk͉�MkT�<��V)_��
n�GPl�k�6�5Hc5#���~6mp������D�);���.�����Z��HH�k\�G�����  H��}p0��)�䴧#�P���d ���  .�����B� ��ʥԭ
�h<�r��R+6PD�K��eSB�(� ��r�H�D�6X�("b��& ��Cf� ��r&��*D��r����20c�rq�U��l�@p�u����������vrr��~~�w�I%#|�)������À$  o���H�7ɇ�݌c�1�c�1�c�1�c�1�c�1�c�2͛(*Ef�۰'���Yh.pࡔ'#�^��s�|���D�,��̭��Q��y�'j,a5�������jښI�%�AXޔɣk���6��P�O�h��^n׬\��noQ4�g6\�ߑZb� �)�-��r��$�͇ײ���4)����2x��MZ1��{h��Po���nIiu�W�׵״W3�3�HE*2�} o�EOQ�w [B1S��v��ƛ�ͺpMJں�{�����5^��#`��h#�@�����l{<y��j��Sb)-s�C�Ty�˪J�б
䨏%h\�r �"D�r�˗.A�1�c�1�c�1�c?���1�c�1�c�1�c�3����������"b��&1�1LAD�1LAD�5�#��{rvG{e�P�Oo����ϡ��������`��99���d3�#�C;>���
T�P`���h\�a�+�.hhh(P���
B�Y�;�VFӺ{u1qĩQ� ���0�U�R�d��0Qv�E�\d�˪1�`Ɓ��Td��P<y��%~~8\���99 **?n�S��T��Y���nTT�z��M��i=�֒�6G\�W���.��"I�-i8�ֿ-�s-~l� 7p'�ߋSO��SUbtZE!I��;��@֨�b� #���^�H޴�[�7����i������I0H��@ڐ6��d��M��"j��5o	�����M��6�T�,�	�^�c���蚜m�bk[�&���������Wc�Z$y@�DǑ��P�&����U9I=�Vp��"b��N_;���Q��kM��ʉHx��T���2���k�	V�̭���	jgF�Y@x��%� �+RՑ�4x	��kj�_�jCB�حjN!���Bj�
K�Ȓ4�G*B��m�		5�v�X�$RmT�Sr�i�
k2R�%���C��S8N����>��MGa�Ѡx�vtۗ��$�Z�bUC�;����МD�17��X�ؼ �w�O :E�ݹj���V��$t'�rF�l�H�򅉹�x�� �h.Е)s- �;>���b:$��h9<�p��@b:��#�2erT�.�P��L�A�� ��̜Td�H�?.q+B�K�"�e�X�͔K���r
�.T�L�e�P�2�.A��b��6l���*D��L\� ��r��)�/� )sCC"���b$H.]��B�
������~�$F�]qĥC�i�kZ�kΈ�!���cY�@` �d�ּ�jt<�����c�1�c�1�c�1�c�1�c�1�c�J�y+E��R�2����R�v��v� xa�����sPNS��|�>F��2\�N*G9nx��SӚݭ	iK�6Oȇ��k����wY�$	���$�l���E0H��S���!!4M���T�Ko�J��-�R�W�4����-�:7�2B6y��8���"7~��1���lW�#h�#	
�Ikg-�z���ꀧѳ����~�r(n����'��zT�dQ̭��4|��N#Wk�6�<���`���9�+ow�7d{F�D*W2��v�
�LA
�U!2qQ��4.�x�V���A�b �1��c�1�c�1�c�1����A�c�1�c�1�c�3����������"b��&1�K�D�K�D�K�D�K�D�Ǖ4<(5����2����M��>. 2�%�-�����6��f6��H�$Ol6�������ۭ��`���J0eG�X���2��LX�F�����Q���J��V!))rꋗT������.*9�E˪.]P��4.�ɕ�R��*4dɕ˗_��6` A�&8p�ۚ{t���5!7%0����j7o�T�����p꜑di̹7G_[��	�bk�X��S��F�@iZ�z�\BGu�!ЮH��T��q#�:�#��hz�Nf�%5�a#zy�N��3t�|Kq5�ub�ҳ,���=1�N*Y����.�,��2F��ءP"�T�c`��!M�O�`���~P*_��6������p5�&���S���SQ�H�܉�f���'>���)8��F׬� e#� 4���Dtj�M���Hד���5!�bRtT���h��4�T��a-�1�m�ښ�n�r�~L^�w��ۼ�ֽ�z�\I����mnF�A"4��$N$MF���L&��ȓPE���YS5�%`����:�BJ�A���z�W楘����Z�LF��בdLx�Z@ޟ���A�$Y;=�/�["nY����+)\���A5H5R�5���!$�9~�'��"GAd2م;4 p���hG���G��)�䴧)NQ�*.1�T��r�r꟟���'��
20�����e)�L�h\�rB�6lٳe�4.\��f���er\� ��1�l�b.B��4,\�&�˚����Ô��X��H�.d`���`+�\���~�I#GC;>��U��=�9�G����ϡ��P<�c�1�c�1�c�1�c�1�c�1�c�1�B�&Y.0���OJ	��q�H�%.r� ���VNGX��iX�x���fJy�S�a�x  6�a"5٪}8q�������2p� �O��ޣ�Zi���J���3�$N+8���e�lػ�ȩ0��8:ٽ�T�}T���Al�d�lK��1��`|�|�GLr}F�i��AUP�T�x'y�M�~j�"��5��ֵ����u�(�9 O(>>#i�K^ϔO� ��&w��r޾�Ǣ��X�T4}E�ҠÈ \˓��#�bTT'�T��8�p�A� J�2��)U4.A��X�͖!b!b!b!bA�g�cAH�.\��c�1�c�1�c�3����������"b��&1�K�D�K�D�K�D�K�D����<����tIZ(��R:su����8�*�.�--w��v��p,����{�~nTaeR�O���L���(3����s�z�TqC9�d�a�~T:����%ۦ�Ϯ��0c@�u����%}{2��d2:Ts*�Dd����Ў�y���4.�$p@�ߟ�������1)N*J0�qC=�� ��e�P&���Nw* Y6J��ݏ�Mi0�4S`������h�5M��u��֤4�f�a���+,$'R���YN���OF�BI����$��@�a� 9S�Nϧ����#���Hޟ;�N��j�Z&�K�yM�Mq�@ӡI�),�Si�$iS8�v >�$ �@	0��P�L#p9�GZ�ۮI�״�5�{tMNn$֐7�%�YL�&�T�&��*oI�b@��1�CV�!:
m"Ę�I��d�ى`�R�VAw@�j�&��@׫jl["o_L��HLVV���MH��a�KH�	:ԁ'[Ԭ�7�'[ZF���D�oT��1Xw'��I��|+�j��6֚U�c8�˽��:<��ǫ^���ΰ�jWo�i!9 ��k�9�^������%�8+"knZ��/�(ՑI����bV+�[f�y�L�P�6G�V���o�jWzh��:�F����y���{T��a���D����.)Q���U%�h�h��T������	��A��4��*`�J���Ү\�Ȑe��ʗ*D�6lٳe�4.\��f���er\� ��1�l�b1L�f���0`  p��A�c�� �"D��͛"�A94�C?Y�d� ��ն�L� �HY�c�1�c�1�c�1�c�1�c�1�c�1�l�Jp�S��.A���4)K��B�>L?-7J�^���#��\��3�o���Zi�RA֩ ��{��c��u��0M����H#�{ �O��.Tq��L���HFw6���B��М�e���Zr~j��U���d�� ���S'�����.<�03��g�4F4E�]��Ċͪx�a#��9�d�� ��aB�`3d3�c��}G�s{LOs>l=�'�s��R#*�����ˏ���"���c7�֊�'�_m
���+B8��݃'��fq��IZ,�d�$�Dйr�J�%<���IZ*D�6l��,B�,B�,B�,B�( � �1�c�Ar�˗.c�1�c�1�c�1����c�1�c�1�c�1���("b��& ��Ce�.A�.A�.A��6lЙ~G}Nrsl(>��#�{}ONPL?j�	�:
Ci��޷�n��T��ܨ����ᔮ��͖�e���P�G���)�O����	���14�1�M3v���[n��0򣋌�h2]�X\�ˢ~GT���ʢ�Q.�`Ƅts���21�������;;?4�nG�����������S��>���	��R��B!תa��ۙ�`��ɲ�J��8��L_�J�4�6����Ų2%8���b*RF�D��ɱNLo໩��SC�4BV8
�U�5�;�ՏV��:�!wRh��L$o[#���hz��r�Y�=MGe�I�:���J��Vm�B!�!I��:.v"-y��<cL�l�N��F�r*�H�`�~Hn�I	�,]�dE������S��j��S8^D��4�vz�V cU)���4�V��i��wY���;zI��N�x�GdbsȖ|���N�y�`�)�L�e�jl5��mj��S���y���Wy�%S)(���jt�Ub���;����\�+4�Jp�U�5Y�5]� b&�rד����I���I���J�5���b��SH��+�!I�$ji�]��E��Y�W7@ͮ���l��-���e�!5��Sj"_/���U�Vj��/#���)$K"%�Ь�IKD�N�i]Nm��	����� �0���Tpb#�X�-q�A�9t@�s}�0�Ɔ
.ж�������]*䪘d�"�W%T�2����<�6X��l�D�M�*D�&Y��(h�\� ��1rb6X��D�6l�1R�FL�2d��˘�"D�r�� ��1��1� �"�]\����܏ʋ]��y��.2p���۽Ꞙݴ*�c�1�c�1�c�1�c�1�c�1�c�1��*h]d�s�K�8e('7�ǕY\yU�/��G�F��I_��4.v2�wg�ÚP�6��� �K�I�әhD(�!�*�\]*:۰�a1F��i����k[�Kn��*�'�u�<]1�����LGn�E4Ӈ��fW;�[\�2�	Ó&fL���V��N.��S��3����wr(72D�L~~>vS�� D�x�Bf|�~*PGl�P�:�F�E�D��hc��kd��ZD�,�|�{E�Ch\�v�Dʤ+�Cf�1���"Ar%M
�TйL�f�ٲ�,B�,B�,B�,B�3��� ��"c�1�c�1�c�1��f͛6l�AD�1LAD�1L��("b��& ��CeLAD�1LAD�&1r
��8(`7��17�b�I8�e��94���I&�4�kZ���dT66���L>>G1+B�r�L�<й!߀ �D��� NNj�Q��BO&��6�M&	�:��c =�2��?P���ĳ'(�P~�Qv�s*� . w���oc��  ]���IAG  ���f�u9��[{{p�#ǘy*�����! �I$�I,Z�7��L�~�l�����qjzb5��8�d���1���}>t/�F��=�n�5;	����wA�t�B$k�OR�r�!+��4"I�Vd1��ބ�����e0�$SX�T��yS��t$����Ȥjn]f�3��YnV����ܼ
���U~iz��S���V6��`��LD�q��ٲF����s�U��b�"oJ���nLH<�!@xj�%��@�Q�hD`�)��m�]�i6?��-���)�D�J�á��4O0kJ��r�Ș�}7S����%�(�_�Ʀ
A�9�6��y�����m�l��j;-	n#��l!�)����jX����tx��&�T�1�F�cx6�&����#��5��h&�
e�ԍoMּ�iY���mב��~Z�+@r4ЉdLQ����Y	8J�w����V+�MD��Lm�l��i�C��@��,F�͑$�Ck�ԦY��3*��q���G\\R�/�E%8�y(ƃ#�eC;.� at��.�hb��''����.y�B9���Wh@a����ˌ2�&YD�2͔K�Tйr�H"e�,B����1r\� �L��A.AL�f�:�˗.\�3�D�$]$_��%J�=�������>#7#sl�����G�e��q�11� J	�l��1�c�1�c�1�c�1�c�1�c�1�c��2͑@�4.���Bxa�w��_��#�2�ʀd�e܏��9?WW2��`��yHw6������"I��ZK1�J�	��~6F)���k�ש�4�����P\�
d�R:�'8����6��GF qu�Nm���NI��A���s&L�.p3�ڠ�Z˿7_[mTO��;NnM�g����"�����(�B� 4/E��о�9��S�`#܎[��K#�`�ʥ�M�b$E�]�˞h\�,�"����OG��0�뛙�&P��aB�����=�8qr��Cf͖!b,B�,B�,B�,B�?��c�1�c�1�c�1�cf͛6lٲ�r� �r� �r� �r�!e�PD�1LA����& ��"b��& ��"e����jM����#T����H��}vn���������{{Jp�'��7dL�<x�,�2��Ў��`��I�K�@����~�w�[���t�g�No�"І �R��\�D S@G 
8����3��ggg� ��20RS#  .p�!B����	���(;d ��a� (0�h�iA�d�@��DN��`��ǝ��QS����`ȬT�5	7�'֪��6�nｵcp��M�s�4�t	���.�Y�ƓZѯ�܊��o$�&���VmA�����|ډ��iS�JU���T�&�M��\��ip��b�A5�Y5�MGe�eL֓����۸KRF��Q&��|D�,�/�������ރJ�g[ZBQ	5�t�5�6j66\R��VZ����`�)
F%�0�V)	����t����nG%Mkr�S��D�R�D�4� ��0u�M� ���<wl��.�[��n_�	��L�:ޝ���E
By#^ܵ�'��0�N:7/#��8��>z�J��	dЬmDMぽ	&�Sc���OF�#�JN!�A��t!<N������㠚܏�FH7}����S>)�����#����i�l��S`9�j��&��^Q����% �Hj�|�v>X�)�#hI�&�2<`�w��M<ħ%�"��(W糏��{TP�[s(b�@'9�} 1ʢ�Q*BЊyt�BҮ\�FC?G�0q���.B��H�.B͔K�Tйr�H"e�,B����1r\� �L��
%�.T��,ٲ�&1�T�R�J��v1���"D�&1��"hJ�bަ�%#TL�����IE#�{ |PT�t,���P4���8'�$,�2r�1�c�1�c�1�c�1�c�1�c�1�c.ASB�'�D�#��2�^͓/�� ?eq��+��*OL 0l��� q��mP��ƃ��=��O Y:�꜑�$�6�� �|�s7L �P*z�?n�*�%A����2�%�:�O�i�e��.��:Tp��h.e�=@��xb9�����=f���� �Q��l��ng�9#�M���6�YH�M	 >J���s�Z�
��([�����`�5P��m���4�	�c� )-*��Y��m9�SB��P�" ��e�3� No���Y���r&��3�������b!�f��H�%h�f��T�SB�K�bK�b,Cf͖�ʬ�Uf�q�PD��Z,��R�����8z��H�#�h<�ʦ��Ud��*����4tm��i�.]�Hh\�Р��Jd��g��Wx�~�����ᔦK���r���8�..(�gg$�w#����Ѧ�I����e��t��%8�P���%GG<)��2:QE�̪]���˓��ۘ��a��K����)�����GJ\bS'8� ���fC
h1q��R���q��`���3�@���;fZ�Q⢅�8$���2$��^]@u*ف,آ1�I�-���햫��$ڄ�����$�D�&��!�|� e��98�W�	��YjinA�PjM�:��#�ڃ]Q��e�p6�e�cꀚ�M�bpV�ፗzH��tԥK`�ZhO6�7��rw6,�M�qk��#��\�4�����֓�Pk��w6	6�%���P�%�
N!#Q�q�1��	/�A�֭p�CSr�l��RD��J`�	>o��2Ț�/ͭɴ����d"t�k���m4R_���mx�8��F���ۤ�Ԑ]��eD�Tן�;'�Ee�Mjb	/��CU!�ֿoDJF�vX<J��O�^�s�?9&	�MD�q�`ۡ��;@�u����R��`���k�򵡱\�nڶ�&����1�@ސ�F��8	mWyY+��W!�#[(�QЖ�k�����y�phh2qPaM��9��}q���a�KoĄ���r:9�J�"	��sLLO2eq�+�D�*	R�p�#&W2�ɕʕQ!T�d��Z4 �(2�
V�G44.D��44Lb&1��D�"c1���Lb&1��D�"c1�cD�1Lb!b6X��X��X��X��A;;6S���=�hJ�Q����̌�H�������c�1�c�1�c�<yrT�$H�"T�U�5�
 ����l��D`��i�*�\]���ub�n��Nv���J�~�P(-(w��}}�����  �&`&�P#7�l9�;�S�4�v"S��#c���4UB2�;�3Bے'��\�\��h�d3�����4*\��D�"�e�IZ(C9=�	��H�.Gčܔ�h���D�m萢	��C>�9���<(��a9+�Ŷ��۰#��48p2;�۰�'�B��40���a�քT6�C~{�p�׳�R���)l���ˏ*�eH��
������6X�͛(� �yP'ױ���D�6l�
%�"\�ٳf͛6C ~A,���X���Ǘ.\� ��A#�<��͑����`�Q˂s}Oi�9�92��8q��l>70R7ɢ�2&���a��G1�0��e���)s�
@�Aw��j�xaǷ6����H@�:I�'�IО�s21�`��4.�P����2��q�a���@
8��d ���ҿ#�G�S�B8���9=�s ��SB��d�s�=8z���O���G�K!1�C��U��q���T��B�7�M0���_�ӊ�f	!G�Z�a��I�O$�EFS��ަבܮ�I�ƕ3�MdRY�d�#i�`���'���k2��w��M1"��ZD��	�&<�$��#^&�)�)
Oi�a�#ï#I�5�{L1f�c�dRi �X�:��k��D&���oBJ�Z�r�)4��I\&���Z�!5#��ZOA؈�LH��b6�\6��+��m��#^�mLM��dBV�M�JJRX"3Q!�f|�)(�ޤ�y��tVN��R�����Шj�F�4��kI�1ԑY�wn^Gv���Ml#ME��jqA��ؓ����x��4��
C��)+�̑�Bj���'��h�B6-I�-�h�R�<nq�9��4���f�8������P(Y��*L�NIR�:�񍑳�#iܮ�F��DK�շZ<�N#��5 H�b��4jyi�<ף���f�(��pǞ�4 ���x f���bND1� �?~~8��)98È�D�*�0��%J�È�D��hh�]A
�BЩ��T�Щ��.<�r�H"e��D�"c1���Lb&1��D�"c1���Lb&1LAD�!b!�e�X��X��X��X��D�����C����b$H�A�����1�c�1�c�1�c*T\��)R�D��%˗"D�͛6O#�i��^�u�zi6�D��(?K���ȩ1ȩ1���)�R���GCZ֣�(.������'��ڲP#7l�D����Pw�չ;=M�A�"I*��z4�HK)�7?�8�t���cB�5�1�uR$M�Ӝ�\��4.AR&����5H�8xQv%Tp����"[X�ȓ�i�E
���C��W���\�FAP7?{NsPLl�~GTe+�s�t����PJ R�PG2� P�g��R���..�񔪒�2��l�J\�A��\��&Q2�
&��������l��6X�r�NKno��*h]f͖!A,�
��r� �R%ʑ*h]e�0�ʑY\�8��`�4T�*TH��A!���q��,��a1@�:Z�B�ٳg�"D�R��K� {8\c�r{e0�`�愧<1��'�ң�cd����pge��T���u -�KI�I&��S!A�`j�f�>LG~8���w�42��:9�&W8����v{G[v�P ��^̆ �0c(��{0Ï�N#�h<�̴"�]<�d�Ҡdʁi5�i���GO@��ۑkt���58ӊGB������f�q��|�~(�a~$mNoO��!5�u�����4�\m�;5���Y�)����؉4yA�|�%�5��C�]�Hwl#MDjB`�e��kZ�R��|"7;����jBZqRH�p�Ĭ�;+�C�ԦT�H�ȑ�M4F�����rյ+���RȄHm+�M+7"F�8��;��&�����j�n�P mZ���"$Ґ��(M���[e�Nl�D��4��摴8	�¥!<��4<��W��`�w���Ǜ�Ȝ�oZeN�06�I�w#oO�T��ӣU$K"o�I�f�ND���ND�� m�H��:R$�c��WF��ț}A�G�}�sOj�ft�A6
r�GS�]�iL�OH���H+F��a0��I���A%pU�Wé󇛤��b�X���~iF��I"��dMi%�E��F�tx�]��j�MJr�]�&����e���� R'����%9��?{{��� r��2�����裇8�*Ta��J��8���8���K�PeN%\��S!CCh\�+B�H�CD�"c1���Lb&1��D�"c1���Lb&1��AD�1�X��l�b!b!b!b!��J�ɓ+�.A?A"D�&1�����c�1�c�1�c�3��D��c*T�r�Ǖ4<�+E	��ܛ)��eA��� r]	�R�d�	s��
d�y�?F��)��;G8���~6&H�y����kzWH$[�c���n@����榴�~�ToE<�
ЉQ����Y�cAs�\��IZi����z
� ���Jp��4(h2 Pa5�֙�Fʡ�����-�����)�Eݟ���h~��O~[v vO[.Q�A��~�(0G[v�PO0>vLi��-��T���4P٢b�ʑ4.h8yRV�"2�^��4Lb�,١<e/�������,Cf͛("b%�"\����N8e*S��.B���r� �&.T���ʑY����s�K�2~|��Ll����1�� ��J�*D�6_�
��e��{��{���wd���'dw���J�\`�G#�%K\�� �b� ٲ� ��i� ��(�{MA�A=�A��>0[l�L�V������%����,ךI�i���S���
Ty�L�~ \�uIR�\����0cB9�B��GJ��db�9��{d0c#���h\�8�#�\�ds���2Ў1+��f��A"I4:�o��
� 7T�My��4w'����݋Oѭ��W#X��RE'a3�v��b%h�Zh0X��&�M{��bIbBu)�J&��%�B/"�n�@ڿ�����4�RV5�%r`񤑾'��	1Ր���O"o^Gsc��+�7�'{Z$R��aS�jb;:�@ҧ,m�	�D�y=��$�Hֶ@�%�B��$Hm+���d��sF��'�,�My]�n�!
7R<�iJ��D�'����&���S�[�k�N"u��υ(D:׬�m���jq� Ԙ鵹;��y=�ׄ��󹱵!$CU��4L7$o�9W���Su�Mdn�',�5J�6mP 6�	�xH�H��S��bm���`6j2�&��$�|�u#���l��8�2��w��q��:��27���m�*;`uID�\�H�0_�^Gsa�D;$r�IDWHIͻ�����~�Y��H�5��sxm���B�ZW'��s��&�,������h>R ���*�*<���(R��#�\erR���S��C2\��ts�����8��uFL�8qÈ�Dp�#&W.�`Ƅts�48��S�D)��'�H�4 ��йV�K�b&1��D�"c1���Lb&1��D�"c1���Lb��& ��B�,Cf�����
�ˑ"E�::9���5�$$${{{0b�˿c�$H�����c�1�c�1�c���cA4)K�h8z��������a�9�����eҊNs�h�J`<<D�_�5L�c�Q��kg��~8y���S��2(�`��֓q:�e�Q#�n�i��7���.r�ʑ%h��T�q�TL�1����X�)�ǒ�*J�xa�B$FOr} D�G"PhP���\���2��S�l9�s�2=e�#q�4k�y@�����Z6:�M)�'9�������[@R��T��PL*7��D�p ~sNrLj��s}AR+6l�r�P١J\��������!AD�6l��("a�)Q�2\�%�Y\����"e�(�!f�8��E��UM�*D����R%�q�=������44*T��,�.p�9u�a�~���9ȡFF@H|TZ�Z`|TZ`FD&H�7"l�=��}vTd�#�R��~{sJ����ގ(cA�A� G �]����t��~�7$t(����`�kM%���R�0Ϯ�U"U21�3����%J�È�.���vv~v{G~y*���s*�.0�K�d����G}G��01qO���� ?
 0�FK�80��gài�����T�F�F�����k�B%+ů')Q j�sl�L䶼.�X��N�J�ҥmMo!�x�!+���FշkMcŗ-�n��m6<I���5Z�6�e�I�_��fк�biq��N��L<�4	GV%'2��0H��'$SE&�bSm�D�ju,�-M�)$$�〲kmB�đYJ:�)	���j�N��4��wRȤ�	��EKa#^OD�N 1<�i�Mj�I��F�k��KH�]敁��D�Q�#Sr�R�e5�h��'Z�ЌI�mz̔ީ��U��f��]敀�zo��Q㠈M�i06��	O-����0ꑰ�4�T�V���$w4)ƪS�����������PJMR%��x��`�Q��r֒�p����Q��r��ލN�ԑ��y�{>�"r}*X�[F�W�c�=|�wO$MD6�x�;N6\&��V&���|"0,�����.)�$�̍�Hm-S��΀�ב���wpB�&�(f4*2\��d�4#�@�v��s&W%J�T�
���S�����ĩPGG<��x`Ƃ��.�`Ƅts��矟��d��&W
G8�(�8ĦN*rs{~e�r%�1�r%H�CCD�&Q2��L�e(�D�&Q2��L�e(�AD�1�X��l�b!b!b!b!D���r�

����2d�$H�c�%˗����c�1�c�1�c�? T��T��*[�c��b*�J�(��@\1U+)X�Ɔ��Q9<�2ۓ�z�r�GC�Id��<1m=�&&�(0�N}LOP*?l��9K��<P�p6�k�a>� 7Zd��r�f_��Pٳe���6l�D�,B�S���l�O� ~8(e�)r���M�LU��*[a��R����yA��� ?'�
Nsl�[�S���;=���i��Q��{dL��=�@���`|Alc�����Cz�)���&�H&:DH<6����(�ع6l���ʘ�4-������A*D�R&!�f͛6PD�ʑ.T�͛(� �6R�<�朞��A�DDbo'B��0�("e�K�0b���bbc���T�W.\�&Yh8z��U�mZ����׳�!�EĚ{ ��Pn��D��e	���v�gg3��� {{r[$$_�'��;9�h\�& ��kB:!�� ��H���l�/ڨא���n�%G)��)R�T����~ \�uE˪GG<�TP���{~2 Q�ᇀ
8��������b:�
J01��e˿J0�S���<�\�::9�&UJ�b8�e���Wf����Ф�&��F�B���,��m�5��mI������wmѩ��9"����;���Y�(�j�Hu��MM�L^ZCR�"vF�z�Z���%sȦ�S�����p[r�nJ$RH�D�4�M�L-w�Sț���^&�&5]�b�$�:I��ܽK*cQ�|֐�OV���kJ��5"�$Y}-R�N��R��b5���$ЉD�&���mׂ(Y#Z�|_�T��gst�H�۵]S�Ly�;J��X��|�ce�M7�`$VH:Nj��t�bf�)S^�j���Cf�Gb#h��T�&$���J;d�|)�@� k��6���&����-1�bF��%���F�&���E6ۤK&��m�,�$;�7�NQ�������k׃p|�V��j����4KY��*֪�Ҷ�k�,�d����-��q���1�M�kI�E
E����6ڷ���ȩdel�u$K;��@gA�U~�Z�l�6�"k�bMX)�i#J�f����d�m�`��#�~Tp��Y��
Jx�h~~8(RR��
���3e��(RTts�4�0c@����
J(RS�44O`��<Щ�2d��*D��K��J�\ɔ��*\��L�e(�D�&Q2��L�e(�D�&Q2�& ��"c�ٲ�,B�,B�,B�,B��Љ&1��"hhhT�S���"\�r!�����1�c�1�c�1�1qĶl� �R�X�.Jp��f��T�l�\]��IP8�v��4.�"Nn�[%��:�kpnˬD==� ��@'�˪A��'ӏ�����('��#i0�|6�l��9�=[�"��oO�M̿#�8x�[6l�2͔K�Tк͗���W!f����I��S��2�@e9�
l�%s{*w��E%;j֨5O��~rs��]�����	��.��Zn��i���["eNg��f�a��,�D�h��~H<6�y;� ~A%h��&K�D�1r�G��*h\�,B��w�������\�A�M�"\�ٲ�yR%�Y�e�lٲ�6l�TPZ6@H&DQeA��6@H�S�.q�L�8��A9mm9�ᔨ"b���.]�[i���������_�9�>����~���i�99��mmͲ�~rr �����si����jYi��#��Tx���F@>�=��18��NY_���Ԑ������st�Q���JqQ��	P8]P�IFh{{���\��B����0���cMl���|�Ol'>����00c"�.�pȤ�U"<�S��%hJ�*S�%8xc�$��L��~t����ShHҦu��$��5X��D��֚
�˱���5mք�Y�L95���@MDZ�S<�I2r�kMd3���jR�K+ �դM�hֵLFޚ�z��HBs(o���Ta��:�m{d��`���1j��F�������m�;8	�Kb�Գt ·bE 5<M�{?S�楙�.�tT��B����t���"YjH��%��΂se�ir:,I�WAM=tmJ��1k~7�l���DҺ��4:�N��Ku7� q3����		�p3A֬���F�`�<S:ڧ�\�[��	�E	��d��4���"6��~�;�0w�N"Gn�9:���$܄�ӈȞ��ɽ)�)�Ӈg��r'��L�Z8D�'`G�g���c�HKq	�ɇ��h�|M!w2F��b�:�NoH�Dő9"�)�T�#��J5$BR��@���k&������֐�S��W�L�T��K"Y��I�R
�{^M7 _�6O�;8e��Y��
~h))����S��>��.]R�S�;;?&&'��\��&W2�ɕ�L�.]P���GG<p�&���THPePeZ".q+�8ǰ��a���?"e(�D�&Q2��L�e(�D�&Q2��L���"b��,B�6l������*Tx��˗�� �$H�����1�c�1�c�1�e��ya���HY�D���"Ef��4 �
���/���Uf�
$�K��{��ܛ����ʏG��h�Z��3�2�3����ވP�B�&�HH�y'�=T��17d��w��\p�,�r�*D�1r�Vl�����@�-���M�e���V�=K]�׷�������yN��8�&�> n��%y��;���dL��̥�9G.��O �Ol	�D�Ϗ�2��Pn���R
�6[�3�R�JЎ(e�("cA�H� �R#�Z%hD�!D�������1r�G��JйR&!�e�l�bK�\�%�1
%�*h]fʦ������z�q����ϓ#�~)��P<��SB���]SB�6O%h<p��%<0�As(���T�����t��I�z�#GS����Ǉ��zS�Ǉ�ĝ��"i�o[R�0"F� c�2�c�d3`�R����z`�kS�s����bN��屈��E.�y�*�"21���a� ��̈́��N`�7[H�#�3t�0���#�T0c@�I_�~�� aw�!�?0���N#�.��<��xHjX���Г��lz�[����&��Tѡ�|�!,HN�A-"�@x�$RpZC��1�VQ,N�y]ZI�5�I�6iiF�r[��6#����'��J�jE�L_�]5(IX���K%�"�I`Js?X�l���ٵ)+�A$�6�bSZ��J' �`ބ��"cx�!$�z��� 5N ��.�mDK�4���R0z�K��mj���RL4�6���ƚ��Ԑ�WLz��5)���;�`m�]=t5�'e�c�����kA����X����{�4"^,N��˩�	-��h�k�~17!��\�%���&���Pש�[�y��w���[x"QLJe�Hjܻ�&�漄�$o�6���$�18�����[��Є)<u�8��N��P�{n��i�W�h]sٹ���E!-��������p�%Kk�j�	��GCCzOQ�i6�D�j�'�SJh���3I��R�J��g��8�$el�1��3fq9�m�A� gx"��-�tM��#IIl����4(�����;?�1���\��x �8qL�\p�$�P<y��1*TDd��@��G���A�A��WJ�bP�??#�.q*V�IZ"e(�D�&Q2��L�e(�D�&Q2��L���"b��,B�6l�����T��gA?�`����1$_���c�1�c�1�c����~�p:=��\��*^p�S�Z"D���B)Ƅ2yt���.Dd��ʑY�DybQH��������V�y���g����s(V��%����r�nt�-�"�����Ҁs}}Nr<0�+�b�,�h8ySB�6U4.Jp�8aC�ݓ��ۭ5���^� F�2P�$T�6n��A~�i�GQ�)�B�ܑb� �i�&L��*I&����Hn:FP<�Zn��i���#��Йv�0����P� $��ϩ��˚��z�s�!���4.b1r�G��(6�ܝ��
Jp��f͖1�c�1�c�1�c���"D�$H �Ω�r�H�*D�r"cٲ�R#�Z�ʦ��"e�6VӜ�����2\㳛뛓��K� ���l9�;*h]eLCC<�q���*A?��d��6Q.<��)��ɺ���Zn��n�Q��蘛�a�<�S���YܜBkJd��4��Y7��  ��w�f�H�%2)�����TH�:��������X�	�˧i��ڥghT�' �"hJ�BT�\(RW������������  (���n���
G2�R�]��S��g  �����pS�8  >��~}J)���ydw&5��15�^7ķ�j�L_�O�D% I�t6#	n���MZ��w�b���+7^�Ӎ���H��)��V�u�5���̔۾���8o���3J��b1,�D��y���WsY[F�7�"ȉX�,�&��ޚ+��	�n�a|OtT�#J�̉�P18	� ���[16]�yM�:�����"�����+$K^D�� 5�ښ�SD��$�-I�&8�·��k�Ұ:��b���loA���\���Mi�����1��lMb��Mr�L���+,�𒸩$"R��U�H��+7/;�"����D�$�I�"P�S)����L�k��չV�JkT��5"�n*8�#;$	F f� 3i��8���k����@�ӈڣ�{dud�Z�l���(�!���k��BI����ҍX�MAv��OWl�������V��pt��J��vp�)	��ju99J�)�.e�Ĥt'(�Ғ�$jY�n��@�/���@���qՉe��9	�ʖ-y=DP�)����Y��Z�{OO�ebR�ZE2\�T�P~~8��(P���PB�tɕʕPB�tɕ%GG<d��Phh�.��uH2�'�Jys-
�R9�cu����hm�T�+B�)O8��ĥ�%2��B�J� ��44443��"CCCD�&Q2��L�e(�D��1�c�1�c�1�b �1�c������������" ��f��"\��H!���d���Ѓb�� ��"e�
�(��\ÉO?
�2ۓ�a:�U���B���`��?
\0���L8�͓��@96T����-#kK&�2A�!�m�(�4=B���\P��R�<�RV���A�P��>~7vw��DGD�LH�l��1�eP �2��������	���R��o���gB���l+��K$�s�A�O4
svri��D��� ��\ᔫ�"�f���R'�#�Jp�%�Y�e�X�1�c�1�c�1�c;�Ar�˗.D�΂&1��6lٳf�A�M�"\��)DȊM�����O?>LTк��H�� ���,CeLCCD��1�M	R؂8��Zݝ���zžL*"~NN(L""j�Q�n�y@��tLM����dޯ��Q L�L���z��h���{Mвk��GAЬP�M�M�ԑC��Y�I�����*8Ё�����9 NPv��d��˩R���qAA���`Ë��@Qv��� � (�9�A�Ҁ ]��`g����~.�S����ݓݖ��T�i8��<O�Т!��ŪĘ�z���#BsԚ��@YR��
;j�x
7R(����I�H�:ޚ��d�ݹV��o�j��6<�J�"�)�K�,O��i�$&�!7�p6ԮZ�1 n��4��J@�hґ74��T�Ո]~jY�/�eJr;Ub�6wkN�7�58�<iR��g�����,�^Gv�NVH��SZH��)���ⓨD�(�S���~MA�lQ�bKi����5Z݆ک"�|N;�@�&�i�Բ�wkI�ks�|�t���CԲܕ�h�r��R]I�D��̬���'�|NWM��������R0t��u)Zl|�lG��Aw2$kȲT@֨8�����^�@�T�h}*8�D:��I�ܮ�M	��gp�H�<�*�hړ��5�j)�H����l�b��u�!,Jk[�1J9�˽�5�M��h5�b;Gb�44��ʘ��ik� my��H��#:	jU�YLZ�6��;�$�%2�h$ֈ��	ѧE!1jY+�BH�mN`H�-F�[r\yP���#�hT�K�"~~81�&W2�0c �#� \P��42�*TD��q��3a��d����;;?9��2qR�UȨ2Щ�2�\�S)O!�A��\�"AR$"ArCCCh\�R$2������!����e(h�D�&Q2��L�e,c�1�c�1�c�1� ��1�c?��������=�[l��SӒ���E�%�"\��H.A����$*�� ��1�4 ��1rAD�"b�(��D�Sˆ. 0�g�e6���.�ʦ%T�����>�d���ݟU#��e��ɲ�BĪ�9>�*�&�eD"x4�K�JEf�A��#��4.T����惇�g!� ]���srr$-D�)���f�\�u���<ѱ��}�0�����7��u9���((p8

�J��Ss"��Jq)�1��CCCCC\�"AR$2������1�c�1�c�1�c� ��"\�r�˗.\�1��lٳf͛)NJp��<����}{#"70j�y+Brz��T��!���rS��.B͔1LT��(h"b��ǎ20a�O�E?>�6�i���k�dtR6�#�2D�"!�:��޷��q9�4�O���ڥ�QѲ�0DV��
w֚cL���<�nP�n�P+ '&�[�H���F������,����H�I��7JqP����<�w㏮a��EЕ*˪˛�g���UʠA����PF_@#�� s#T1�`ϯ��� 	m�=��P�o�A"{xl_<�v��ޅ�Fһ��S< �+T�!���m�5�[�rC�^�`�Fּ��T�y9�<KO +�
��HRu7���Ȥ�16�!���[��pYm��w �`�M��saФ�M�D�&��3a��"o[�����I�68K% I�<VX��E5��Գ(oJ�c�İ0p�!u�5�0p��c���j��	$��%(�u"Ȅ�w�V	��k�j�w�V%hmTφ�LJ*o��	���?H@�rrA��4�6�b&�D�@ڛ����"[�#j@w5��wZȘ�n�������lM�z��sh��H�)$���w!��d�`�OX>
���e��.�x�~-߰�c�
rs�t\��F�Po�����F���1��4�l�0I$������8�H��dX?�RD��w+��5վ�	��@�)��jra���PM�ަ���|BkA��8�J�Z�~�j�K.�ʙ�ڕ����Ҧt��#P5dM;5�#[Z"m�b��Ȗ�1�$�c�x�Z"O*w�)Ѡn���N��K��h\���{{ sǘ0cCe��~~��� � )*T�*U1�AAب����FL�}}����J�U.�������#�G8)�8ĥ̴%<�R�$(2Щ��W"�B�(2�
�T44445�1rD�&Q2��L�e(�D��1�c�1�c�1�b �1�c��������cB�$J���ml`�LD�� ��B�("b�L\��"��BhbA��.A��b��& �!D��*�"2x��'L-?���U	�i��5�Ȅ�����*-*$�=dc�#Q,�F�20�g����w��-s
/hEhEf��Y��������_]�Ob�S����?7_Hگ�����0Sa<��u�DP�c49��'�S
����l�5Z��V� dɂ5���)�;�dJ� ��BTLb���4.Dй�H!�����eR$*\�1�c�1�c�1�c�$H�"D�c�3�6l�b1�.A��K��f͔0���aO���#�\��H��A,�Ty+E�("b���BЩ��JШ�ĥ�.0��<��L8)��LuH֚���MQ�j�$P<�F�����S�ǔ�r�! 

	��
v��N4Ri0�������==�T��*N>-.	>xQǵ�k��;�^M��V1��#bDm�2���Jd⤪��PCCBx�  ���ɓ+�bT�#�T��e������b��'9���rr  s�*<�%�?���1 ��nm��tj��څ��xސ�F���)M#Zhu��IX�+$G�U����I\C�!��ud";��/"��xԥF���)(�V$��'5�*RߌBm�=�9���,� �S�4"Q	����"H)��1$�6\��@M�Kw��b�H��!���|�':��v�$�������(oJ�f�+e�Kj����qB�Dq��|�v:4'���bGu����F�E�;?�Zӳ|p�ׁ�I|�������bm�n�kHک�
rr@�W��m"���1,
�x鵹7X���\e�k�k��-�6G��V%�SS�,t��o�M�Ԓ�LH֑V�ͥƧM���q�kd�4H�')+2E�0�bR1׃ a�����Ǜ�eJDsx��HQ;h��T咺�ҦF��I�rE�!(�V%$�&����c�lQ�tt�m&7��cpz�Mj��bNO#M)�bi"kL�� oHOShIHM5��M����սM�mh��.�#<�&ж&�F�0pQ�@i|Nj��W���6�kĝ�@� @�hh\��B*A	�+������)��NPPv)+������.�R�$S�>��i�܏b�S&W.�Q!.e���H��2�0���1�r&�Ȑ��#��G `g����8�)�M
���#�4*b��K�
�y��*D����4L�e(�D�&Q2��1�c�1�c�1�c�A�c�1��������A<������d`Ƅ�W*Ef͖!A���X�r.A� � ��1LAT����e�
�K�*D��c�;dݺ�z�ڭ�I�D'���MH$��o%���Vl�.d��	�i�TR�!�fʅC�Ïo�KT��w���0O�`��@*2�������4T`�F���
-l-���Ѧ	\�F%}n��O�;GO["z�O���G�����\0��*GG��n::��lvs���)͛6!b!�AH�<�rV�G�.T�L�������er\��1�c�1�c�1�c�1����
��&"\��H�4.Tй�W*Dy+@����`�^�]��� �p�[6Z*Tк͛-�J�f�A�M�Y `ds��G�S�8��s#8q�����F" 7���Ba�`���+LD"�!%������R&��k�����d�2�'6�T{e�TFT@�i��9&�$�B;^j%��ƅ)H�ے��s��:%ʏ���us-�L�Ty��)L��`�ND��<���\�_��-�{~20��A�>�G���	P<q�.���pȧ�f�h�~�'5����I\F�X�z"F��g@�j�&+e��^�*t�C��|n�Z�ԑ9�)$��ZO��#zu���1jJY�Dk^v-X���j�d"_5�w�|^:	�#�ĥp[Ƽ$�kM�Og��Qh�%�H�D!&���1��� .��ML��KN$1,�H���!�׷$I��^u����1"�dj�)+����jP��Г���܊0o�CV�yȚ�aCzW$,��J`2Z�حM�ޓ�'��`bY��w�-")�ID��q������,�\���:c���I�8
���8�d5n\��A��jmyM�t7��P$�ԓzL�r�	��k4�qx6��YL�$o��Knא��"k�1��x�I�DkZh-X�� �-7yM�VY����E
JF�!э1&���S�qZ&�!8�j��Z�4���y���*S�Dԍ�kZ�6����d�h�?" Tyl���I0I�kJD��,�Nw[#t>�/�ѩ)��t��w{tژ�mV$Հ�ĝc캁��5FA
 ��i�S����*hd�BH��K�T p ���2es��g��R��T��2��uFL�<y��K�T0cB$*�Q�%\��W�F^�?%hT�T�rCT��u�S1�S.�B�&N*8�qī��D��#�W8����FN<�y1�4 ���S*�TʦU2��L�e�c�1�c�1�c�1c�1�g���������1�a�ǀ  ���  ǕQ2͚�AA� � � � �"\�%� ��"b�D�1�����<�>7}P[NLi�} db��kr����3t����9��hVک��B�hA6T>�\�02��P��B�a�w0M�'�Y����6�yj�̲�]̍��nӊ3hD�n~�#*�3B	�����BZ� {O>>~rrvi�ڤdi͖�L��윞dS�%M�*hD�s*��� ����b&P���2��L�e(hhlc�1�c�1�c�1��� �$K�D�K�\��H�4.TйSB�ʑG.���&DP6@H�n��ܝ�����
~G�er�J� ���Y\�A�J�*h\���ʐD���z۰��%<��s��vv����m��_�Ch�4�k�N��n6ו��յO77ar�bN���떈�۰���пo��1%�h��4x2y�w6��sU�Z@j'�E#�j5��@n�a�@'%��4T��#'�e h� H��
�ɕ�L�.]P���% (� ��.1pA��]*�]\���Jep��\݀'99�b8��j�+)��A�):��F��&�̐�@ڤ��ShI�$ש��&���ޓ�ަ'���ԡ�MY�F��,��Bcxw+�R��	+�D%c�ĥ1,Г�$NQ,DK��R�֩����eJ��'��`fӲh��I�oV���F����g��#F�Qh�Vd�&��$jR��\O"�Hj6+JjP�r�zcmkr�18�$�Qh�<ڬ�CV��5o��r���*U�IXmS�5���=��&+�U�!��%�����d���rYnA��שe�;���FnVR�Q�i���Kr:;�R{խ��N�h\ج!��(���ce������b��S�)�W~�׃GVB'�M"ڕ�	�����k$kM�m���4mMmi��bY��j��VH���tǑ9���;�O��9Yf�P�7G���Q����MtR-W�5�֩�ew	C�ҔR`���t����7A1�&לr$�l�5�epEL�yӇT���jh�Vm���I��]0m�M�P�;�$�HՑ8�ȡNK&��ŉ�Lޔ�9��}~\�@b�Sݞ�@#�<��U<y��O`�IV��� .d���0cA��A	r�hss��R9�'8�R��J���45�1�r$4A�A�HQ!D��WJ�)�IO"8�q����h\�ؤqFNhT�r#ȐhA��ڦU2��L�eS*�D�&1�c�1�c�1�c�1�c�3���������˕*U�Ç����Ǖ ��+PB� � � � � �("b��& ��B�4*��1*#P�*�6�zP�d�q�BCɣ��4w5B� ��f�M,��	&�$$�qR��mR͢oQ��s��s��oքJ��U"H��=��xQr��<�й������Z3,���n�.���
�%�Qˮ �x 
%Ȑ\���L?<1����a'��bޝ {ٳf͍�ArV.y*&1(hhhhhh�D�&W �L�����c�1�c�1�c�1����\�q�ǎ8�R%ʑ.T��.ALAD�,By+C���ۚ�H��{��	��l>�b6X�b9uM���U4.<��SB�M�%h>n�-� \񓊟�
NO[i�[�3�����j1I�s����kM-�d��1�i���y�11����* ���*���Z&<�Y$��R��;�8�����1"z�X�6����i<��tN?(���ي�8d�ħ�J� ��o���˗T0RQA��e���`�^��>��ss���� `dt���?<1w0B�T�S.�8���brp$��e�7g''!O����59�bw4$�&��j��$L0R�D&��j�;��%6�I4vt5�a�AHy�Nl8���NF���Ee*���y�+�J̍dR?_���@���fP���r[xu��9��ii�T�Ԭ�4���� ��ܫMEw�`��.|��k���U��JJ�/8|�<[�0�l?_� d�5!ءbWn���2ɭ�t'�ͧg����G7Y
0o�%%b���kM�����j�B�c���zf�k�/q�R̡�S)�����Hkb�4V)	�V�܉HL6���p�^">w���E��ZO}j���Ά ������E$v���U~�6���S��@ސ��ԆKLy�~�Y����-�AIXiH�SEw��$�k���7y9�jP&��[�#E�KH,���5&6֚�E2�xC)�IJBb���S���Hy�m����Q��Eƹ$j64 0sn��5�����iѠ �q��diY�BS�-=�t|&�,�{(pJ�"�<��N>pM��Иۛ�Z�b��J� k�OV�.ޔ�d���Imm�������	�����r}} ���1���\�x���e��``�Q��.���IR���\�0cB:9嵷�`���<�1)�er*����йV�H2�
�V�L<Ё�4 y��LhT�K��Z0�B�2qS�s#�J��HD��H*ev��L�eS*�TʦQ2��c�1�c�1�c� �c�1���������� ��T�B�Ș�La�&\���T���# ?2���THPEA
PB����,B�&.E\���8��d į�]�	��e��W#�l�iOP�)0�L�H��DP�n|1=��ڝ &69��	�?i�	�;5[�1=̻�&și���&ʃ@T,B����*��s�A��%s{2��q��c�#/`*�=��	&�QRQ��̌ (3��sA��E?'4�/WC�l��d�#�UJy�*��	U.Еu��]�AL�����A��b&Q2����1�c�1�c�1�c� �cA˗%J��r�
\�r%�"D�Lcg�<x�%�t�1��20aA��� �ڂs"���Ǘ44.<��s�l�\�A�H"b�H��2��� 0�r�@?
NO[?>L?j�S��H�-�Z�kMH��I�0�]��3��4x����0Lt{L���~ob�֚`��m��I�i���M�ǝi�C���,а_-��f�*S�#��6�cd�<���r!�� 1��ࡋ�ˢvv~21��G� w70� 2er��ۓ�'��A��GJ(�@dt�o�T�=��GG<1���M���zs���۳�q@��%C�#�I�	$�'gy��Y�D��I��Y�e��mNRk�n!��4����c��	�
s��MdRmJᚮ��Բ�Hחi�_J�&��iZ�F�����X���'�ޝ����SZܖ��f�h�P��(=t�BgC��5�iX-����z�Rkj;�m	:ަ�ݵ	<MG`wy�"H׷'�a��%$��'yY"wR��
�B�����J�!�Qh�t'��Sb0�ے����j�Z/Ʃ�	��%��R�n���#X�zF��G��zBi �D���tKw�rF�.ޓO#hINY+�N��a���k���iB�����V&b4�OX��Ǒ5J�yH����۬A�6�h�Djm�Ew����p�`d�cUdO0M�Ć�ŗ�حoM����Bh��W�g�������YX&;�bF�(j�A؁Ƞ�nS{Ly�H��Ț��t	MD�p�{�j�f�jd%�Ą�p����x;�����'{Bqk��<��mM
'�ܞ~�mD�E6�4�5�Eu����;��-y0����m1��>Ln�J��O�m�*�qrrp&�a�0c%˪	��P��L�1��T� �+�L�\d��P~~81��P2ep'�@�#�B�u)�G�hT�L��A�2�
�UK�
��ur*�THQ!A�D�R�B�G�.2Щ*�J�T�B<����L�eS*�TʦU2��Lc�1�c�1�c�1c�1�g��������J��r�!��}}}b���j	ϩ�IQ��hk�D�HPB���!f�����U.�Eb���k`�>� s}PLl�[vrl�U. ��9ny����@��ݟZ��d$���{�~ӿr(7*t=h�����@f�c�	Ǟߓ���Tع�Z�2p�Y�3&P0�������M���n��Jr��ja�k��{e���l��?�Î����
i�����D���A�b&1��Ub�X��?���������1��"�PPP???{}}<p�G�{ �Û:$z�4 䡝�[�����m���T��MQ4.TЁ����%.e��DƆ��˗"\� @�m6�iij��������N��4��L�m��ƃ�;(&��ė�k�`���DH�*#�.����w)��b'�H�PH�j��<���֪5��6���RqV_G.��`P:nnnR8aH�#�~GG1Q�O��4  \P��L�J��P.]S��g�p�GJ(�@Ë��.~.�(G��ܓ�4����
~hs)����� �L��P<�-(w���[%�jȈy4w%�My,�md��<��F(A�������K�E� �]���Ul��Z�5L�� 7GP$�j���ӡ����ZF�|l;#�Z�pm[w�ZۭAu�M�;5M��a$"~5)�NZA8l�M5�	C�0�Q����jA�Nw	/��i]������\J��4_�M�Q�D�����	��)4�6�~iY�J�E���f�&��!�Ԛ���G�bWp���]xc	[��Q�j�%5�g��ҰMěV�x�k_�R-�������+L�LI�6�Y͂I�czMq,J�V�e4I�V�A�|h}+:�㢙�w5�����9"�o���E�KQ&�婥1����t�M�"#����RI�E$�Ԛ�J���N_	��A�f�o�J�9
\�\�0x�H�8Jm�HiY���C��Hb��u	i9e�S�Md���&��[/$st�b���r�_!
��Wm�W�C�k��P$��L�yHčo�c��\��&	MQ��BH,I�%+�"����[��CM�@j4�����B졪�n~�{{��y���:9����;?�\���  .1��Phh�2�ɕ�̴*]GG<x�G-*l�����2\���PT��T��%<��B
��
���%<�)�G�T�L�D��H.A��b���Lb&W �H�T�H�h\��r&�Ț"<�sB�K�b&Q2���1rD�&Q2��L�e(�\�2��L������������1h\��r�˚.C\�qÇ�d`���\��,D���AR%ʑ.T���+�b&X������ ��TL�b���? }{��x�UIZ%h2�]0�@�݁'6�֚se��0���I�R��UHO.��T�[`|)��~�* >F���:M�`����s�{MA)s��o�4�j�i�i͂�n��`������6�S%߀=�{{D�RT�X�
)���  D� �$A��D�"cX��V"c����������.\�*UJ�"D��r�nnj

��8e����~ y�.͈1Ƅ���`` �ӗ2�	�9���	*8�/��s.��R�WT���Q?<\�B�LA*Tdɐ@�7[�׷��Ǐ�����4۩��6�g5�
�P6$�oZ����^�srGy��dM�3�C� ��3r�i �d��`:$�oV&�kzb�)^Fּjvo��RE�����M��d��?
 `�B���?#�~.�� � �#� ]�rꋗT(RW��_�
8(���U
2���@t�� ���% ���
�� ��g1H�)�����R�T� �"����dk��Cے`�u��o����黁0MH���S�V��Z�~��r0y6H�/��0M� �Oe��t�s���'����ZZ@(�M�w��M��Z�6+^Fš��`�����d�IX�:jmA�5��4��`^�����%�[�ֽNVY��&��'�����jk1,	E����	0X�	D�E&��Z�&�j��қ��ךd�r���:�n�)��x��
�9IjV5���ZAGoB�4�5 ׄ�m�I�iX�D�Qi��D֝�����jyȡ�F�r0yM媴ZM��m{r�$K7oMo�Rp�M �):��5�zW7�ԋ�ԦM��B����)��M!Cz�tW�"j�1�RF��"j@�N"M���=LQ䴃qmTςCkr�D��	�,��Y�ٵp�����K 6��<����I�����Ĥ�<ڟ=M$���̀NoJJg����j� ���~�*N> O7w�=Z҅9���(,�ѭ�]0��p5���^"')�M��P�sl	�	�GBi�d�P&�˓��Ӝ�#��˛�` �d$p��� \ ﯢ������  ]��``�A=�G�$r��>�0-i�-� ���INU4U4ObT�hA�S!T�y���%<��B
� ��H�T��1r\���Lb&1r\�"AR$"A�r&�Ț"<�sB�K�b&Q2���1rD�&Q2��L�e(�\�2��L������������AH�4.\йsB��hj�*2d��B�ߟ��
J�1��AR%M�4.\�%�.A��\� �!��("c ��K�"A*D\a�O��K�TйSB�("b%� ���"8e)q�OJЕ*�'('-���-j�(N$N$ Pn����Pr7>rn�_[
6��@��� ��As�2�3A��T���8��C����~|윟A�ʏ�.�J�+CCB �444*T��b&1��D�*�U��D�!����������aÇ�*SǏ2e���  � <p��Q߃.��lA��A�߃9��l��\ g�峂���70O?7��(��ʗ*a��
.�0��M"D��J�*PPP_������L�hhhj�Z�I��nA�]��GTe��-p&��Ѩ�)ͦޖImyL��kM+���P�7F�9&��Z�햨��&ɹzm%�A�6��Orj����Ijbr�\K+��kW�ʎ"\��g��a�� ~G)�0����<���8`�_��??{{�����  ���Ҋ.ЎeP�*��� GJ��q���D�৳��0 ��O`��rN?(S�"#I]�l;�ۨ�O��6Qߓ���Tᕷ�2�����~S-1���Jr[��hoHBGB���Op��"q��~6t �w�G������6)	��(Hu�$����Z�2b�dk��/RL���F�ԭ�]x�:jR[���_-:��|��~,S�������h*IJ�$��@��VX&�k^v|�~?t6HEI"i����:ަ5��pMד��|Z�����JwS�K"m�lx�`�Z�cđ�S#N��Q�ބ�$�hk[�k�D�oJ�F��`�)�n�6�睊��rq�$�F��䍫nFjq�Z���X��E5��!ݲYl�S�Z��YĚ'�����p��jLj�măqkBH��.�t��4i�m�R�F�����֭���#:�@ײ��8��H�L_�[L#o�گ%��zMm��y=~֚�m�`u�$o�M1�Բ�V�Z@+UdRLpM���P$�uS!���
�I����4jp꜈�Ow��#�!W1�'y��55�J�#��5.Km�2!��"��j��ݔ�S�D�*���m7'��O��2(RWgg���Ooc�����T���>��i�ݟC'')+��9��a��b8�E�"Jr����x��@�B
��
���%<�)�G�T�L�D��H.A��b�D�"c1��b��*D��H4.DйB�G�.h\�rD�&Q2�.A��D�&Q2��L�e+�b&Q2��444?��������H�4.\йq�J����ǟ� ���*8�M�4.h<���ʕ4.T�H�T��1�X��X���\��"c�h\y+B�H�D�K���R%ʑY��R%ʑYJd͕��� c�gsh���<bmD΋#�Cԍd�r0j��Znm�����G�ʤHT��V�� 