3611
100
100
1
223 1
39 01111
224 011101
48 0111001
37 01110001
46 01110000
195 011011111
241 011011110
123 01101110
133 0110110111
199 01101101101
188 011011011001
69 011011011000
246 011011010
136 011011001
240 011011000
114 0110101111
122 0110101110
132 0110101101
158 01101011001
190 01101011000
251 01101010
115 011010011
135 011010010
218 011010001
238 011010000
214 0110011111
235 0110011110
232 011001110
248 011001101
57 0110011001
59 0110011000
134 0110010111
213 0110010110
144 011001010
208 01100100111
67 01100100110
54 0110010010
34 011001000
202 01100011111
86 011000111101
93 011000111100
68 01100011101
157 011000111001
160 011000111000
204 01100011011
94 011000110101
101 011000110100
108 01100011001
162 011000110001
185 011000110000
118 0110001011
200 01100010101
80 011000101001
83 011000101000
126 0110001001
26 0110001000
23 01100001
247 011000001
43 011000000
221 010111
253 01011011
129 010110101
211 0101101001
142 010110100011
149 010110100010
172 01011010000
111 0101100111
117 0101100110
140 0101100101
210 0101100100
119 01011000
230 010101111
35 010101110
255 0101011011
22 0101011010
29 0101011001
186 01010110001
187 01010110000
226 0101010
131 010100111
193 010100110
50 010100101
177 01010010011
178 01010010010
138 0101001000
254 01010001
47 01010000
40 010011
175 01001011
217 01001010
28 010010011
31 010010010
109 010010001
237 010010000
128 010001111
215 010001110
32 010001101
127 010001100
231 0100010
192 01000011
76 01000010111
170 010000101101
179 010000101100
14 0100001010111
15 0100001010110
85 010000101010
164 01000010100
88 01000010011
103 01000010010
110 01000010001
145 01000010000
30 010000011
173 0100000101
209 0100000100
60 0100000011
206 0100000010
205 010000000
234 001111111
163 001111110
113 00111110
49 00111101
120 00111100
252 0011101
147 00111001111
75 001110011101
77 001110011100
71 00111001101
159 001110011001
165 001110011000
12 00111001011111
153 00111001011110
91 0011100101110
104 001110010110
96 0011100101011
102 0011100101010
183 0011100101001
184 0011100101000
17 0011100100111
81 0011100100110
90 001110010010
196 00111001000
121 001110001
167 001110000
36 0011011
116 00110101
139 0011010011
191 00110100101
61 00110100100
189 0011010001
216 0011010000
41 001100
207 0010111
4 00101101111111
10 00101101111110
84 0010110111110
99 001011011110
20 00101101110
212 0010110110
233 001011010
38 00101100
194 00101011
219 00101010
198 0010100111
156 00101001101
171 00101001100
79 00101001011
146 00101001010
21 0010100100
51 001010001
201 0010100001
181 001010000011
16 001010000010
78 00101000000
52 001001111
55 001001110
228 00100110
244 00100101
250 00100100
243 0010001
225 0010000
45 0001111
227 0001110
42 00011011
249 00011010
53 000110011
130 000110010
242 00011000
245 00010111
137 000101101
56 000101100
229 00010101
58 0001010011
166 00010100101
169 00010100100
64 0001010001
92 00010100001
98 00010100000
125 00010011
72 000100101111
73 000100101110
66 00010010110
100 00010010101
105 00010010100
151 00010010011
152 00010010010
87 00010010001
89 00010010000
95 000100011111
97 000100011110
70 00010001110
107 00010001101
143 00010001100
106 000100010111
148 000100010110
150 000100010101
154 000100010100
197 0001000100
25 0001000011
155 00010000101
161 00010000100
236 000100000
222 00001
220 0000011
33 00000101
27 000001001
24 0000010001
203 0000010000
44 00000011
74 00000010111
174 000000101101
176 000000101100
82 00000010101
180 000000101001
182 000000101000
112 0000001001
18 000000100011
19 000000100010
65 00000010000
168 000000011
239 000000010
124 000000001
62 00000000011
63 00000000010
141 0000000000
vinicius$Qj[o-�"���H4t�ӧN�:t�ӧN�:t�ӧN�:t�ӧN�:t�ӧN�:t�ӧN�:t�SSSSSQӧN�:����u�����������S4�El궭�QQQ[f��:�)րhj
������������������������������������������������������������������ւ�j�KRhQ,+kd����m[:Ԣ��[:S�P��$
X�V�XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXA)4I$�I�U�(�7ږ�Ɩ�TIV���Na�KM�&��G�<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x���I��Lpd�A\�cB��H�th�D�l���8��M5H�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�07 4��qq"��F�X'N�4�i'(b�ı\
�i��i��i��i��i��i��i��i��i��i��i��i��i��i��i��i�be�.%���$�oI��V��+lձs����TqR�LA��������������������������������������������������������������������45\�R@�Fف�5c�cKgI�5h����Ѡ�)�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�M4�VNp�7��(��e�z6�6���,h�֑H�\�=�{����{����{����{����{����{����{����{���x)<��5 ����֥!\[����PqTt��#�6bl���{����{����{����{����{����{����{����{��)c�!\�H54TZI�L��X�0ڹ$JPI9F���{����{����{����{����{����{����{����{���d��@�Q"�t���N��9,d&�	[č�[��7 W��{����{����{����{����{����{����{����{�����'"�[%%Qo9���SVX��QL"yc��^���{����{����{����{����{����{����{����{�c��'�P�Y屡��yEl
���pF�2CME0Cr
a=�{����{����{����{����{����{����{����{����l��lC$Q55V����Th"��cP�+Cco6����{����{����{����{����{����{����{����{��ǘ	p�E�Β��	p=Lڲ6�Ɔ��������{����{����{����{����{����{����{����{�
�<�m��4��	F��I�0���Y!��:)�AJ&a�a�a�a�a�a�a�a�a�a�a�a�a�a�a�a�a�a�i#P��P�Za�a��)�:��X
� m������������������������������������������������������������������������
�-����d��������������:V����{����{����{����{����{����{����{����{����{�����Ě�\�,'=�{����5!`)�c��&�i��i��i��i��i��i��i��i��i��i��i��i��i��i��i��i��i��i�6Qd2
&ͦ�i��i����!�����{����{����{����{����{����{����{����{����{������1�{����.[�i���͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳf͛6lٳfޭ66b��f͛6lٰUh4��jT{���������������������������������������������������������������������������*�X�c����������X���Ph�����.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˗.\�r�˭ �N8 ��.\�r�˥1SED��L�]u�]u�]u�]u�]u�]u�YraR�"
����Ra�*TB�S9QDːHw]t�]u�]u�]u�]u�]u�]uЅhi�L�]u�]u�]u�]u�]u�]u�]&DLϱ�D+�u�HD�Jg�f}�-�ˇ��u�]u�]u�]u�]u�]u�BM�k`�9�뮺뮺뮺뮺뮺��
8�T T�4*�3��M��L��������뮺뮺뮺뮺뮺뮺�
!vh�9���eK�&]dZJ�͆�3>��>P���oG:�]^�\!�����%f�	���v����Z)EN�
��6��Ƨ5�'������
kl*h�.�B�뮻��Q�7����v���Ҋ���,
  l�V�X8�R`��H��%��]u�
�����BDI�����뮺뮺뮺뮺�(Y��E�� �ia�f��3��
DB:u�Cu�]u�]u�]u�]u�]uۡ
"V��00ru�B�]u�]�u�]-��+NA�� �qqL@���y�s!5 4��O ����]u�]�뮺뮺�Ѕ*�`s�����W***p���H��A��JB���=��ż�X��xni���t��
�=�(ֽ(�Q��*Q~Lh!B�!B��[� +�*���T�W�s��clz�R���Clu"˚m�jʏG�֣&��e�+;3) #d3��Q��t�q29)r�!B�!Bҝj[H4M a *�뮺뮺뮺�@�<[I���nM�+B��YV��N#%�����c�& 5�mx�l�VI�X�`�m�@R�Uҗh��뮺뮺뮺룂9�l�� ��*T�R�J�*T�R�J��+�@�r�N-Ǭzסƹ�k&�>9^J.�g�@�C�)Mr�۲�x6��	��
.�Z+��U�J�*T�R�J�*T�PG
�-�ƃ���뮺뮺뮺�D���J�4�
��I�n��"�RV�	��o6��Rm&�dā$�� �&�!JAD�eEK��뮺뮺뮺����Y��3�N�����+�\%J���̔$	b� 	5$���"g7������+i��3T[���Y��4.��eJ
s�"�몆�뮺뮺뮺���v��P��>P�( �@d읓�Hch	i[1��)JS�i5�0�:HJ�hm6����N�3��(��kh�1Z�1���&�bQRZVE�@  �@  -6	��4��S)��e2�L�S)��e2�M!$R���$O,B� 2(6�i��h3F���ie��3��DF	"�`ŀE�+dLX�"��n���A��e2�L�S)��e2�L�S(M- b�kFH�cZ&&&&&&&&[�+%���cR�i��&�H�`�"40�l4*<��8��r�#����Q`�Qh:�L���M�@��3��X��-����������������N�e#�M`�ģ��j1�F#��c�F#��l[��pF�dx���N���	h�!��g�07C ؗ*#DZ�g�-bч:��碅&� �)��u:�N�S���u:�N�S�,l��mXG��M�n˲�n۶�.�kFMke��G���D@F�f���5.44"!&i�d���0�L�9 e3�3�+e��� Հ�6�r�nF5����j�Z�V�U��j�Z�V�V��9�Ȕ-p��ŷ77777776�hũ��<�I& ����U���h+�M��� b�)<f��G���6�m��Q�`R��P�LlY�q�&&&&&&&&&&&&&&&&�nB���h�5�����q8�N'��eĜVf\�p�9ۭRG�rjR{��=��+,ˁ�^sX``�H�SRQ �K�Q�+2m@��2<<nnnnnnnnnnnnnnnnk�,����b�B�&���*
���*
pc ,RB�U���ň�� �m �Q4�E����Hf��'��M�$Qi�Q��HCRD��TM��kP��an8�5$��`0��`0��b
r��Si�h���Eu�T�Jh�%Q˲��,��3l��=�]S4�B���͌�"ǋ	�%dې4&���H�*�0Őh`��0)�p+�-:뮺뮺뮺뮺PH0J�ZKd�|!]p�lA�*�2d�E$%T��}��$g�$�(�,��ћ$z�1��[T�W�b�@܁V�9�D�iD�q*�=V\CD0`��0`����i� �jmc�	YYYYYYY[}Lh���YI8�95S�$��ymfMM˗.\�r��fQ�E�P�Q�MG$!��R�Ԉ���Jl�����Z�NVVVVVVVVVVVVVVVV"7�i)!iX��3|�L�S)��e2����&�YBı	�
,J�[[A����.\�r�˖eA�x�:0�?�����&���`
O,�Hę�ةN�S)��e2�L�S)��e2�Lr��iX���iM���������S��bh�Q"	qBjB�o6�N.4�9˗.\�r�J��#������*
�"Y�
,�x��Y�2�+%��l5��YYYYYYYYYYYYYYYZ�L"3Y�D�k
d3E��o�����}��T�����X �۳�����E�\�r�˗(�`��m(�[��ɊPI�qp9�i1���7ҷ����}��o�����}��o��D��.��b�ehm���������h��l`�k��F�����g�J c5{�.\�r�˒�@sV�jg��0e�`y@h�4	DU� �@�4E*X4T͆�1�P��s�����������B�X+A�M7�1��R����`��r�˗.\�
Mķ��LX6�=f^�N���+im�Vs���CCCCCCCCCCCCCCCC�\\�S��!l� E˗.\�r읓�(R�ʲ�ڃ.�Ki�QYPf�A@f�˗.\�r�̚F��3�c$� n&Ԥ��i��:)V�a�T�.\�r�˗.\�r�ˬ��Fhк�L�뮺뮺誢ЅM��Nl�-�$��#&Ҋ��+�.\�r�ˁDXmJOx�́����Eh(��	T�\  `���u�]u�]u�]u�]�TH�A뎪T�R�J����Lbm��:�k���Fp%�q1�R�r�˗.\�r�˗.\�r�˗.\��@j-�� H�LM$˅R�J�*T�R�J�*T�^�Jf�.$�g��0p8���)P�LK�t���jq9C4\@��qf'��r�˗.\�r�˗.\�r�˗.I��꼉�b�)�������p8���p8e

A���BHHE��H�R)�E"��egi�"��6����%1��g-���p4��˗.\�r�˗.\�r�˗.\�r�X�4�ػR�kQ�M��B��E"�H�R)�E"�H�R)ײ��'i�X�b����������`���BN�i�!6��3� ���É9˗.\�r�˗.\�r�˗.\�r�\a��m�e��lxŞ5�{. g���7!SSSSSSSS湋<c%��,q8��<@E 4T��zz��˗.\�r�˗.\�r�˗.\�r�#����LZƃ�qp��SSSSSSSSSSSSSSSTy�H�A�Zbk��������4cp��Ųes ��]�l0ID�c�1a�\�r�˗.\�r�˗.\�r�˗, h�����6bA"�nnnnnnnnnnnnnnnnY�q2`��O�)-�����������"�,7t�M��`��b���'�r�˗.\�r�˗.\�r�˗.\�6�	��V&��=4k2�	�������������������!V�ܤ *ѱ-��e��l�[*u�LZ�B�� f J��	������ܹr�˗.\�r�˗.\�r�˗.NqD��D��8WL�FC&�e��l�[-��e��l�[-���Z&�u���JJJJJJJJt�*T@��N0J��ң���c��P�(�\�� ��rzzz3=F�����}����(�`T��Qr�����������������P�(��
�H:8p�Ç�W�"TZJ�k�4�@5��*� %9�3���c0̏PPr������DK f�lƚ@�a��RL���*�s$�g �8p�Ç8p�Ý*h�d���"�Ŏ�����~?�d�$�e�� �`��F�A�h(���L��'{0���˓���L���h]Q#`]֒�"=$b4SAJh�?������~?������~�h�9[M"j�>>>>>>>>>�5gk�v,P��lR�Y�i�S��v>OF�3׼AʕAA˗'���j��"R(+���Fs�4�Y�R�BT�	$V��B��P������������� $��c�*�9S)�Y�@L��!�0=Ȗ�j
\�===X�.
�Q�V��h %U��(���կXXXXXXXXXXXXXXXX8����0�YϚ�5�����������G�Ow��D6`F2�F���R�m�zl����.OOOY �Ba:E�]�iYZ�$�Pe�V@�-�U�aaaaaaaaaaaaaaaa�nmȍ7��-f<k��6�M��i��ky����B,H�1�,,���(�o��*�(���.OOO@�$��	(	�!Z��	$�6XɍX��i��m6�M��i��m6�M�|׷$���qk�".��5�.�)Ř�mz�Z�6�����%h&jje�G:3LPPr�����M4�M��к �62�2 ���P����,�6�ReZ�
@ �i4�M&�I���E��h�Z-S��5'�� ԫ:<d"���+<�[j
,�3��rG�P����l6�� &�Y�B��W'��2���L����i4�M&�I��i4�M&�I�-m��h�a���.��R�J�*T8p�ÇL�-,�9I
-r=	h ���@��QQ[:4Զ�H�0N��IDCM�Rsl�a�m�"�.�g�*T�R�J�*T�R�J�,����s8��W]u�]u�]u�]u�q2��,�i=�1��)Mp�"�f�����H���(�x@�D�%:LpbO�z�$�D�g+�����u�]u�]u�]u�\@:thh�ZTϓ"8p�Ç8p�Çh�T�gٖC��(�6�!�� �#��h0H�[L�A�JM�kM65'&�d�cm�Vs>^�Ԁ�Ç8p�Ç8qA���#,hª��]u�]u�]u�]qUyS<9�d�' 0T�xi���5�����%`�Y��-�
aŉm�hLl��̫$㔓 ��T9)*�뮺뮺뮺�9�5��J ��%_�B�]����#8�Ҝ�$!��ͼH)A�b���MV,mA�&�
�V�Z׬�j���MZ
 ���g"W�������	 �S�f���!B�뮸0`ҋM,�8�h���M�. lB�NzʌX5X8�X�z=ģ�b�
�!�9�� h3��@#�
��!B�!Z%Aj^q0��t�>�-���q��l0�y�WD�FM��H L���nY��K&�6�x���\�4Y��-%%.�@� @� @Q+S@+����!e�
f=)�3��j�"�92	"P ��&
� ��J[D�* ���!D.��
������T����+��� �,6�F�����k�s�A+,R��^TЫ'���Q�4��a���W�YD�x�!S�0l��^��AAA���WS�\b�S,^*���!D.��
����� *ceD�)a@QV�N	qI�(4�&!� lP�m���tL�E@����(�δ�
����TTT9_h�Y��MJ!Oy� ���e1Ȉ�ui@����b
�.�����
"S� �B����dh�h�T*�,�*	��H"@r��.�4eɕ�[ ��UP�����)րW!\?��]ih�V��iR���.99^Lσ 8�W
P�r!����!DJu��C���v�A^��T@ ����b�R� �]u� ��RaUN�]����Q�6	��]��������]u����u�]u�HQ]��������C���뮺뮺�KB�-�A]����������]u�]uԪA��H�:T��������������]u�]u�a�D�xUpd~����������뮺뮕3�'TV�BK�~������������뮺�3x��ڋP� ������������뮺뮈�Z��V�'�5�����������u�]u�F��3Z�TI�ʕ �!B�!B�!B�!B�!B�!B�!B�!B�!B�!T�p�`ꊊ�Զ���40�]u��4Z)AB�!B�!B�!B�!B�!B�!B�!B�!B�#�Zo0N��jڶ��������H$���Z-"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H����h��ڶ��j�յ�Z�����$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�$H�"D�))))$H�j[[j$Vյm[ 