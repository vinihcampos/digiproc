s���������(++++999999999999999999999999999999999999999999999999===999++999+++((>\�
��
�NNNNNNNNJ������������������������






















w˝��s�������������������w;���s�������������������������������������������������(((((((((((((((((((((((++++++++��(++++===99+++5555=9(�������������������������������������������g3���s>[�g3���|���g3���s9��w;���s���r���32���������u��s9��r����������������3333333333333335eeeeeeeeeeeeeeeg''''''''''''''''������������������������������������������������355eeg'''''''''''''''''''''''''''''''''''''''''''''''''����'%eg'''%eeef��֧�'''''''%eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee�'��"�3333333333333332��������33333332��������333333333333333333333335eeeeeeeeeg'''����''%f�����%2��������33333332������������������������;���s���v���s����;���s���w;���s���w;��RRfffRRRRRRRR�s9��w9IIIIIIIIII��������������������������������������������������������������������������������������������������������������������III����������������������������������������������������������������ӓ�����������kkKSҲ���������������������������������������������������������������iis�(((((((((((((((������������������������(((((((((((((((((((((((((((((((++++++++++++++++++++++++++++++++++999===<<<<==99554�<9(�������������������������������������������w;���s���&fe.w3���s���w9IIIIIIIK��RRRfffRRRRRRRR�s�����������������������(((((((((((((((++++++++++++++++++++++++++++++++99999999========================<<<<<<<<55555555555555555555�����((((+++99999999999========================================<<<==999999=====+(�+==999999999999999999999999999999999++++++++++++++++++++++++=<(7[�J














fffffffffffffffj































��������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNOOOOOMM-MMOM---OJ�j






fffffffffffffffffffffffffffffffe%%%%%%%%%&j
e%%%%%%%%%%%%%%%%%%%%%&fj
fffffffffffj


�fffffffffffffffj















����������������NNNNNNNNNNNNNNNNNNNNNNNOOOOOOOOOMMMMMMMMMMMMMMMMMMMMMMMMMMMFffj


������NNOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOMOOONNNOOOMMNFfnOOOOOOOOONNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNJ�������ͥ*��-�































��������







����������������NNNNNNNNNNNNNNNNNNNNNNNOOOOOOOOOOOOOOOOOMM----��---MMM----OJ�
��������






fffffffffffffffffffffffffffffffffj
��fffffffffe%%%%%%%%%&ffj

ffffffffj


����fffffffj















��������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNOOOOOOOOOOOOOOOOO--------MMMMMMMMMMMMMMMMMMMFfj


������NOOOOOOOOOOOOMOOONOOOM--���OONFoOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOONNNNNNNNNNNNNNNNJ��������֡����²�����������������������������������������������������������������������������������������������SSSSSSSSKKKkkj����kkkKKKKkkKSҲ�������������������������������������������������������������������������I�����������������������������������������������������������������������������������������������������������������������KKKKKKKKKKKKKKKKKKKKKKKKKKKI����������������������������������������������������������������SSS����ӓ���KkjɢKS�SKћ�������������������������������ӓ�����������������������������ά���������������������������������������䬬����������������������������������������������������������������ڲ�����в�������������������䠠��������������������������������������Rf����fR��������fffffffffff�������������ff����������������������������������������������������������������������������������������������������������������������������������f���������������������������������������������������������������������������ڲВ�R�zmjrxxxxxxxxzzzzzzzzzzzzzzzzzzzzzzzzrrrrrrrrrrrrrrrrrrrrrrrrrPVzzVPrVVVVVVVVVVVVVVVVrrrrrrrrVVVVVVVVrrrrrrrrVVVVVVVVzzzzzzzzzzzzzzzzzzzzzzzzxxxxxxxxxxxxxxxxiiiiiiiiYYYYYYYYYYYYhh__hhhYYYmmmmmmjxrVrrrrrrrrVVVVVVVVPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPP)3PPPP3)PPPPPPPP33333333333PPPVVPPPPPPPP333PPPVVPPPPPPPPVVVVVVVVVVVVVVVVzzzzzzzzrrrrrrrrrrrrrrrrzzzzzzzzzzzzzzzzxxxxxxxxxxxxxxxxjjjjjjjjjjjjjjjjmmmmmmmmiiiiiiiiiiiiiiiiiiiiVVVVrrrzzzrziIEkjjjjjjjjVjYiiYjVjjjjjjjjjjjjjjjjjjjjjjjjxiheehixjjjjjjjjxxxxxxxxxxxxxxxxjjjjjjjjzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrzzxxxxxxxxxxxxxxxxxxxzxxxjjjiiiiimmmYimmmYYYYYYhh____eeeeeeeehhhhhhhhUhmiYhYmrjjrrjjrrrrrrrrrVVVVVVVVrrrrrrrrVVVVVVVVrrrrrrrr33PVrzxxPPPPPPPP33333333PPPPPPPPPPPPPPPPVVVVVVVVrrrrrrrrVVVVVVVV9UmzVVrxrrrrrrrrxxxxxxxxxxxxxxxxzzzzxxjjiiiiiiiijjimmijjjjjjjjjjiiiiiiiiiiiiiiiiiiimmmYYmmmmmmmmhhhhhhhhmmmmVVVrrrzzzzzrzY9@jjjjjjjjrjijjijrjjjjjjjjiiiiiiiijjjjjjjjxjY__YjxjjjjjjjjxxxxxxxxxxxxxxxxjjjjjjjjzzzzzzzzxxxxxxxxxxxxxxxxxxxxxxxxzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrzzxxxxxxxxxxxxjjjjjjjjxxxjjiiiiimmmYYYmmYYYhhhhh___eeeUUUUUUUU________<l_mijzPPzxVrjizrrrrrrrrrrrrrrrrrrrrrrrrVVVVVVVVrrrrrrrrVVVrrrzzPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPVVVVVVVVrrrrrrrrrrrrrrrrU_irVVzxzzzzzzzzxxxxxxxxxxxxxxxxzzzxxjjjiiiiiiiimmYhhYmmjjjjjjjjiiiiiiiimmmmmmmmiimmmYYYYYYYYYYYhhhhhhhhYYYYVVVrrzzzrxxzrrjYjjjjjjjjjjjxxjjjjjjjjjjjiiiiiiiijjjjjjjjzjmYYmjzjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzxxjjjjjjjjjjjjjjjjjjjjjjiiimmmYYYhhhhhhhh__eeeeeeUUUIIIIIIIIIeeeeeeee<l_mijzPPxxVriizzzzzzzzzrrrrrrrrzzzzzzzzVVVVVVVVrrrrrrrrzzzrrVVVVVVVVVVVPPPPPPPPVVVVVVVVVVVVVVVVVVVVVVVVrrrrrrrrrrrrrrrrYixrVrxjzzzzzzzzjjjjjjjjjjjjjjjjxxxxjjjiiiiiiiiiYh_ee_hYiiiiiiiiiiiiiiiimmmmmmmmmmmmYYhhYYYYYYYY________hhhhVrrrzzzzVzjjzVrziiiiiiiimjxjjxjmiiiiiiiiiiiiiiiiiiiiiiiixjimmijxiiiiiiiijjjjjjjjjjjjjjjjiiiiiiiijjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzxxxjjjiijjjjjjjjiiiiiiiiiiimmYYYhhh__eeeeeeeUUUIUIIIlll9llllllllUUUUUUUUUhmiYhYmmhhjxiirzzzzzzzzzzzzzzzzzzzzzzzzrrrrrrrrrrrrrrrrjjxzrVPPrrrrrrrrVVVVVVVVrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrzzzzzzzzxzrrrzjixxxxxxxxjjjjjjjjjjjjjjjjxxjjiiiimmmmmmmmYh____hYmmmmmmmmmmmmmmmmYYYYYYYYmYYYhhh_hhhhhhhh________eeeerrrzzzxx3rimixxjiiiiiiiihxxhhxxhiiiiiiiimmmmmmmmiiiiiiiijjjiijjjiiiiiiiijjjjjjjjjjjjjjjjiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxzzzzzzzzzzzzzzzzxxxxxxxxxxxxxxxxxjjjiiimiiiiiiiimmmmmmmmmmYYYhhheeeeUUUIIIIIll99l999WWWXWWWWWWWWllllllllIeYYh__YlX9himjVxxxxxxxxxxxxxxxxzzzzzzzzzzzzzzzzzzzzzzzzjjxzrVVPrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrzzzzzzzzxxxxxxxxrrrrzxjijjjjjjjjjjjjjjjjiiiiiiiijjiiimmmYYYYYYYYimYhhYmimmmmmmmmYYYYYYYYhhhhhhhhYYhhh___________eeeeeeeeIIIIrrzzzxxxPzmYmiYhiiiiiiiihxillixhiiiiiiiimmmmmmmmiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxjjjjjjjjxxxxxxxxxxxxxxxxjjjjjjjjjjjjjjjjjjiimmmmmmmmmmmmYYYYYYYYYhhh____UUIIIlll9999WWWXWXXX<<<<XXXXXXXXWWWWWWWW4<Ie_hixWDW_mYjVjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxzzzzzzzzxxxzzzrrzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzxxxxxxxxzzzxjjjjiiiiiiiiiiiiiiiimmmmmmmmiiimmYYYhhhhhhhhimYYYYmiYYYYYYYYhhhhhhhhhhhhhhhhhhh__eeeeeeeeeeeUUUUUUUUIIIIrzzzxxxjximmjjmhmmmmmmmmhxY@@YxhmmmmmmmmmmmmmmmmmmmmmmmmYmiiiimYmmmmmmmmiiiiiiiiiiiiiiiimmmmmmmmmmmmmmmmjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjiiiiiiiixxxxxxxxxxxxxxxxiiiiiiiiiiiiiiiiiiimmmYYYYYYYYYYYYYYYYYYhh___eeeIIlll999WWWXX<<<<<<DDD@@DDDDDDDDXXXXXXXXg@9IU_YielIYmhYxiiiiiiiijjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxrzzzxxxjxxxxxxxxzzzzzzzzxxxxxxxxxxxxxxxxzzzzzzzzxxxxxxxxjjjjjjjjxjjiijxxiiiiiiiiiiiiiiiiYYYYYYYYimmmYYYhhhhhhhhhYYh__hYYhhhhhhhhhhhhhhhh____________eeUUeeeeeeeeIIIIIIIIIIIIzzzzxxjjmYYjzrxmmmmmmmmmYz_EE_zYmmmmmmmmmmmmmmmmmmmmmmmmhYmiimYhmmmmmmmmiiiiiiiiiiiiiiiimmmmmmmmmmmmmmmmiiiiiiiiiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjiiiiiiiixxxxxxxxxxxxxxxxiiiiiiiiiiiiiiiiiimmmYYYYYYYYYYYYYYYYYYY___eeeUUlll999WWXXX<<<DDDDDD@@44DDDDDDDDXXXXXXXX<9IUl9lIxYYjjhhiiiiiiiiijjjjjjjjxxxxxxxxjjjjjjjjxxxxxxxxVrrzxjiixxxxxxxxzzzzzzzzxxxxxxxxxxxxxxxxzzzzzzzzxxxxxxxxjjjjjjjjiimmmjxzmmmmmmmmiiiiiiiiYYYYYYYYmmmYYYhh__________eUUe__hhhhhhhh___________________eeUUUUUUUUUUUIIIIIIIIIIIIxxjjiiiimmmmmmmmmmmmmmmmmmmmmmmmiimmYYhhYYYYYYYYYYYYYYYYYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmjjjjxxxziiiiiiiizmmxjYhiiiiiiiiimmmmmmmmmmmmmmmmiiiiiiiimmmmmmmmmmmmmmmmiiiiiiiiYYYYYYYYhhYYmmmimmmYYhhhUUIl99WWDD<<<XXXDDD@@44444444444GGGGGGGGG44@DD<<WW99lIUU___hhhYY_YmmYhmjiiiiiiiijjjjjjjjjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxjjjjjjjjxxxxxxxxiiiiiiiijjjjjjjjiiiiiiiiijxjmYmimmmYYhhhhhhhhhhhhhhhhhhh__eeeUUUIIUUee__________UUUUUUUUIIllIehYh__eUIIlllllllllllllllllllllxjjjiiimmmmmmmmmmmmmmmmmmmmmmmmmYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmiiiijjxxiiiiiiiixmYjjhhiiiiiiiiimmmmmmmmmmmmmmmmiiiiiiiimmmmmmmmmmmmmmmmmmmmmmmmhhhhhhhhhhhYYYmmYYYhhh__IIll9WWXDDDD<<<<@@@444GG44444444GGGGGGGGGGG4@DD<XWW9llIIee___hhh_YmmYhmjiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjxxxxxxxxxxxxxxxxxxxxxxxxiiiiiiiijjjjjjjjiiiiiiiijjjjjjjjiiiiiiiihmimh_hYmmYYhhhh________hhhhhhhh_eeeUUUIhhhhhhhheeeeeeeeUUUUUUUUlIUUI9X<lll9WWXX99999999lllllllllllljjjiiimmmmmmmmmmYYYYYYYYYYYYYYYYeee_hYYmYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYmmmmmmmmYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmYYmmmiiiiiiiiiiijhhjjhhiiiiiiiiimmmmmmmmmmmmmmmmiiiiiiiimmmmmmmmmmmmmmmmmmmmmmmmhhhhhhhhhhhhhhhhhh__eeeell99WX<<@@@@@@@D44GGGgggggggggggggggggggEggG4@@D<<XW99llUUeee____Ymmhhmjiiiiiiiiiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjiiiiiiiijjjjjjjjiiiiiiiiiiiiiiiiiiiiiiii_hYheUe_YYYhh___________________eeeUUIIIhh__eUIIeeeeeeeeIIIIIIII9999lIUU99WWWXXX99999999999999999999jjiiimmmmmmmmmmmYYYYYYYYYYYYYYYYlIUe_YmmhhhhhhhhhhhhhhhhhhhhhhhhYYYYYYYYYYYYYYYYmmmmmmmmYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmhhhhYYmmmmmmmmmmm__iihhimmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmYYYYYYYYhhhhhhhh______eeeeUUUIII9WWX<DD@44444GGGggEEEAAAAAAAAAAAAAAAAAAAAAEggG44@DD<XWW9IIIIUUUeehYY__Yimmmmmmmmmmmmmmmmmmmmmmmmiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjiiiiiiiiiiiiiiiimmmmmmmmmmmmmmmmmmmmmmmm_hYheUe_hhh___eeeeeeeeeeeeeeeeeeUUUIIIllUIl9W<DDIIIIIIIIIIIIIIIIhUW<<l_mlllllll9WWWWWWWW999999999999iiiimmmYYYYYYYYYYYYYYYYYYYYYYYYYllIU_hYmhhhhhhhhhhhhhhhhhhhhhhhhYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYY___hhhYYmmmmmmmmhUemmhhimmmmmmmmYYYYYYYYYYYYYYYYmmmmmmmmYYYYYYYYYYYYYYYYhhhhhhhh__________eeUUIIIIlll999XX<DD@444GGggEEEAABBB77777777777777777777BBAEEgg44@DD<XX999llIIIIeh_eU_YYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmiiiiiiiiiiiiiiiiiiiiiiiimmmmmmmmmmmmmmmmYYYYYYYYmmmmmmmmYYYYYYYYhYmY_e_hh___eeeUUUUUUUUUIIIIIIIIIIIIll99IIlWX<D@llllllllllllllllll9WX<D@WWW99999XXXXXXXXWWWWWWWWWWWWiiimmYYYYYYYYYYYhhhhhhhhhhhhhhhhIUUe_hhYhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhYYYYYYYYhhhhhhhhYYYYYYYYYYYYYYYYYYYYYYYY___hhhYYYYYYYYYY_IUYm_hiYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYhhhhhhhh_________eeUIll999WWWXXXDDD@4GGgGGgEABB777766666666666677BAEEgGG4@DDDXWWW99999IeUIlU_________YYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmYYYYYYYYhhhhhhhhYYYYYYYYhhhhhhhhhYmY_e_h__eeUUUUIIIIIIIIllllllllIlll9999eUUIll999999999999999999(���2��3�   """,,,,,,,,,,,,4��������44444444444444444444444/��������������������������������4444444444444444444444444444444444444444444444444444444/��44,������������$�,��4���������444444444444444,��������444444444444444/�����������������������,,,""  #������������//5�///////������������! �����  ,,,+����6+��*���������444444444444444,��������������������������������������������������������444444444444444444444442��/�����������������������������66�������������������������������U[���[[[VVVVZVZ��YW�������������������������VVVVVVVVVVVUN[W�VVVVVVVVZVVVVVVVZ��������YYYYYYYYYURNU���QQY��P�͆���ח������������ח���������͍�А�QQY���NV�RRRRRRRZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV[[[[[[[[VVVVVVVVW����������������UYU[[YYUUURRRRRRRRRRRNNNNNNNN[NU������N[�����������������U���VVVZ����������������������������������RYV[VZ���������UYVZ[VZ[VZ[YYYYYYYW�������������������������������������������������R[UZYYYUUURRYUR[U����PPP���͍�ח����XXMMMMMMMMR��������׆�͍А�QQY�����RRUUUUUUYYW����������W���ZZ���W���������UUYW�������������������������YYYYYYYUUURR[R[NNNNNNNNNN[NNU�������������������VVVZ����������������������������������W�YW��[YYYYYYYYYW����RNU�YYYYYYYW����������������������������������������YYYYYYYW�R[UW�YUUURRRUUR[�����PPP���͍�ך����XLXXXXXXXMMMR�����׆����АQQY���N[RRRRUUUYYYYYYYYYYYYYYW����YYYYYYYYYYW������������������������YYYYYYYYYYYYYYYYYYYYYYYUURR[NU��NNNNNNNNNNU�����������VVZ������������������������������������������VYUURNOYYYYYYYRW�ZNRW���������YW���R[������������������������������������������������YYYYYYYW����������������������������������������YYYYYYYYUR[RYW�UUURR[R[U������QPP���͆�ך����MXLN'���q8�N#SSSST������cct$VvtsDDDDDDC�Ņ�s��������Ĕ��UUT��������UVVVU��������������VVUUVVVVVVVVVVVVVVVVUVU����UVVVVVVVVVVVVVVVVVVVVVVVVUUUUUUUUT����Ó���Ó��uuuuuuuuuus�uuu�������������������Ņ�������DDDDDDDD����������������VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV�T������VVVVVVVVƆ��tC����������ĖU���VU������������������������������������������������VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVUUT������T�����Ö�Õs�DtttvvtTT$#sa�����SV���d2�C!��d�����������!!��yxl���		��� ��aa]]\����山�%%%��������%%%UU��������������UU%%%%%%%%%%%UUUUUUUU%U}��}U%UUUUUUUU%%%%%%%%%%%%%%%%%%%%%%%%������]\���]]aaaaaaaaaaa]]aa`��������������������������� �������� �����������ѡ��}}}��}}}}}}}}��������������������������������%�]�U�U�UUUUUUUT�}��]]�}}}}}}}}�%U�}}}�}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}������������������������������������������������UUUUUUUU%%%%%��]%%�������]\� �ѝ�����myy��! Յ����?�'�D�Q(�J%�D�q8�Y�A���00a55Hokk^66BBAEEgGGGG444@@@<<<XXWWWWWW999llWWWWWWWWlllIIIUUIIIIIIIIUUIIIllllllllllllllllllllIUUUUIlIIIIIIIIllllllllllllllll99999999l999WWWXWWWXXX<<XXXXXXXXXXX<<DDDDDDDDDDDDDDDDDDD@@@@@@@@4444444444444444GGGGGGGG44444444GGGGGGGG4444hh___eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeel9W9U_eUUUUUUUUUleh_lWleeeeeeeeelIU___eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeUUUUUUUUlIIII9X<lll99WWWWX<D@4GgEEEAABBB66^^koo55a0q8���C �Q?��b!�D"�B1�~?J%C ��00aaHHook^677BAEEEggGGG444DDD<<<XXXXXWWW99WWWWWWWW9999lllIllllllllIlll999999999999WWWWWWWWl9WXXW9lllllllll9999999999999999WWWWWWWW99WWXXXXXXXX<<<D<<<<<<<<<<<DDD@@DDDDDDDD@@@@@@@@4444444444444444GGGGGGGGggggggggGGGGGGGGgggggggg4444hh__eeeeeeeeeeeeUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUeUlIUeUlUUUUUUUUIIUUUeeeeeeeeeeeUUe__eUIeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUlIIUIW<@9999WWXXX<D@4GggAAABBB77^kooHH000q���D�Q?��@�|>�����|�D"��c����?��F����mk�cf��HH((����������������
�������������''-��'''''''-��''*�����������	'(���)''''''''*����������������
�������������������������������������������������������������������������������������쬬�����������������������������������������������+
����������)+�-쬬���������쪩-���������������������������������������������������������������������������������������������������������-���*膇''*��������((HF������mm���'��q8�J'�����@�P(
�A��|�D"�'� ��q8�XMR�����͍А�QQQY����������������NNNNNNNNNNNNNU�����������U�PM�U������������������������������������������������������������������������������YYYYYYYUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQQVNQ�RRRRRRRRUUUUUUUUUUUUUUUU[RUUUUYYYYYYYYUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUR[�RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR[N[NNU�����QPQQPP���ך���LN'��q(���b |>��-�p�7-�rܷ-�rܾ/��
��`�|�F(�Y�C ��a5HHokk^6677BBAEggGGGG444@@@@@DDD<<X99XDDWIXXXXXXXXXXXXXXXXXXXXXXXXWWWXXX<<<<<<<<<<<<<<<<<<<<<<<<<<XXXXXXXXXXXXXXXXXXX<<DDDDDDDDDDDDDDDDDDDDDDDDDDDGGGGGGGG44444444GGGGGGGG4GGGggggAAAAAAAAAAAAAAAA67AEGGGGEEEggGGGggggggggGGGGeeeeeeeeUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU7k4I<liYIIIIIIIIUUUUUUUUUUUUUUUUllIIUUUUeeeeeeeeUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUIIUIlWXDIIIIIIIIllllllllllllllllllllllllIIIll9999999WWWX<<<DDD@@44GgEEAABB76^kooooH5a0q���A��F"���n[��fٶm�fٶm�n��~_�
ȇ���qd�F&���k��f����H((������憆�����������������������
����������������������������������������������������������������������������������������訨(((((((((((((((&��(����訨�����������������쬬��������������)))))))))))))))))))))))))))))))-��,�������������)))))))*����������)*��������������������������������������������)))))))))))))))))))-�+�)))))))-����������������������������''*�*�����������訨(HF�k�m���	�.#�!�q8�O�`�|��-�p�`�Y�p�'	�p�'4��lۂ�7��
����D�q?��XR�ח��͍�АPQQY����������������������������������QQQPPPPPPPPPPPPPPPPM��QY����PPQQY���QQQQQQQY����UUUUUUUUUUUUUUURRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRPW�V^UUUUUUUURRRRRRRRUUUUUUUU[RUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUURRRRRRRRRRRRRRRR[R[U�NU��������PP�����ך��MXMXLG�AĢ~?����~[���f٦d�8J��(J��(O���fY�X-�n���ȄC���qd�F����k��cf���H((����������憈��������������������������������������������������������������������������������������������������訨�(((HHHHHHHHHHHHHHHF��(�訨(HH(((���((((((((������������)))))))))))))))))))))))))))))))))))))))-����ꪪ������)))))))))))))))-��)*������������)))))))))))))))))))))))))))))))))))))))))))))))'-��)-�*퍍������'''''''''''''''''''''''''*�����������������((F������k����#�Ģ~?����n[�f���"Ȱ�=C��=C҄�>�e�f��[6�������B1���?��XMMR��ח��͍А�PQQY�����������������������������������QQQQQQQY��������QQPPPP������������������АQQPPP�А��PPQP��������PPPRRRRRRRRRRRRRRRR[�YN\A񴔔�������������Ĕ��������Ĕ�UUUT��������������������������������������������������������s�Ĕ�Ó��������Ó�����������������������uuu�����DDDCCDtvvvtTTT$#sa���a���V��q(���G��~[������(H���FH�#$d���2@�="Ȳ��8Ne�f���n[�P|�F?N,�T�������cctTTVtVvvttttsDCFtSC�CCCCCCCDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDCDtttttttttttvvvvvvvvvvvvvvvvvvvvvvvvtTTTTTTTTTTTTTTTT$#st$$$$$$$$$$$$$$$#t$#sssst$$$$$$$$$$$$$$������������������������������������������������C�E��sc��������������������������Ĕ�UUUT��������������������������������������������������������uv�Ė�Ó��������������������������������u������DCCDtvvvtTT#ssa���涶�V!�q(���@�rܷ6f����"����31>'����|O��f,œ2G��C���8Y�h͸-��
���E��00a55Hookk^6BBBAAEEEEEEgggGGA4@AooE9444444444444444444444444@@@@44GGGGGGGGGGGGGGGGGGGGGGGGGG4444444444444444444GGGggggggggggggggggggggggggggEEEEEEEEAAAAAAAAEEEEEEEEAABBB7777777777777777777BBAAAB7666777BBB77777777BBBBIIIIIIIIllllllllllllllllllllllllllllllllllllllll@jYX_eWU99999999llllllllllllllllllIIUUUUIIIIIIIIllllllllllllllllllllllllllllllllllllllllllllllllXW9lIIl999999999WWWWWWWWWWWWWWWWWWWWWWWWXXX<<<DD@@44GGGGgEEEAAAB7766^kkHH5aq��AĢ~#��pY�[4̜$Y�H�Y��#�x��<G��(%��b�Y3&(O���f�lۂ�� ���~(���#ST�����ᱴ$$$$TTTTVvvtq�sA�C ݱ���������������� �������������������������������			��������������������		��������	������������%%%%%%%%%%%%%%%%%%%%%%%%T�� �]�������������������������]]`��a]]��������%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%����������������������������������������]]]]]]]]]]]]]]]]]]]]]]]\���� �����		�������my����!���00?�J%���-�r�3l��E����2fbpJ	#�x��8G�#�p��>PN&d���>�>�i�n���|C��!���?�0�����7���������! ������������������������������ #���!#������������������������������������������������#�������������������������������������!!!!!!!!!!!!!!!!!!!���������������������������������������66666666666666666666666*�," +�66666666������������������,,,+��666666666666666666666666666666666666666666666666666666666666666��������������������������������,,,,,,,,,,,,,,,""    #������������!������5���$0��F�D�F����n[2}�����PH�>G��H�"�T��R*E_�_���|N&dτ=(Ne�p\�|AA�!D��?��MXMR�׆͆��͍���А��PPQQQQQQY���������������������PPP�����������������QQQQQQQPPQQY��������������������Ѝ���Y���������QQQQQQQPPPPPPPPP�����������������������������͍������������������������͍�������������������RU�[NNNNNNNNNNNNNNNNNNNNNNN[U����[NNNNNNN[NNNNNNNNNNNNNNNNNNNNNNNU��������������������������������QPPPM���͍���ח���ML����Q?���Źnl�d[�d�ď��<|���0��8�8�8�8��	|�G��8,Œ�	�p�ٷ�~_P|�Q8��#T��ᱱ���cccssst$$$TVvvvvvvvvvvvvvvvvvvsCDvtT&vvvvvvvtTTTTTTTTTTVvvtTTTTTTTVvvvvvvvtvt#cctTTTTTTTTT$$$$$$$$$$$$$$$$$$$$$$$$$$#ssccccccccccccccccccccccccccccccccccccccccccccccf������������������������T��uus�Ó�������uuuuuuuuuuuuuuut�Õus�ē�����������������������������������������������Ó���������������uuuuuuuuuuuuuuuu����������������DDDDDDDDDDDDDDDDDDCCCDttvvvtTTTTT$#scca���涶��SV!�?�O�@�)�n[�m�f���|,���<G���0���A�A�A�A����	|�#�x��L�e2̂ٶ��|ADc�D��?��XR�ח����͍������А�����PPQQQY��������QQQQQQQQ����QPPY��������PPPPPPPPPPPPPPPPPPQQQY��PPPPPPPQQQQQQQQY�P���АPPPPPPPPPPPPPPPPP�������������������������������Ѝ��͍����������������������������������͍�����������NNNNNNNNNNNNNNNNNNNNNNNRR[NNNNNNNNNNNNU����������������[U��[NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNU���������������QPPQPPPP���͍���ח����XLL��D�q?@�ŹpY�[4p�d[�f'ď��8|�����9�@@@@��0�	����>pY3�J��-�����b�Ő?��MR��ח����͍�������ЍА��PPQQQQQQQQQQQQQQQQQY�QQQQPPQQQQQQQQP��������PPPPPPPP��PPQQQP��������PPPPPPPQPP����А��������������������������������������������������͍���͍������������������������������͍�����������NNNNNNNNNNNNNNNNNNNNNNNNNNNNU��������������������������U����[��������NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNU������������������������������QQPPPPPPP��������ח����XXLN#���~(�H����n[�m�fY�,=|,����8|���N�O��������������� Pt| �N�.�/�|���d̐="϶e�n��>"�'C ��0a5Hokk^^^6666777777BBAAAAAAAAAAEEEEEEEEAAAAEEEEAAAAAAAABBBBBBBBBBBBBBBBBBBAAAEEBBBBBBBBBBBBBBBBBBBBB776BBBBBBBB77777777BBBBBBBB77777777666666666666666677666999999999999999999999999WW999W<<WWWWWWWWXXXXXXXXXXXXXXXX9WXXXXW9WWWWWWWW9999999999999999999999999999999999999999WWWWWWWWWWWWWWWWXXXXXXXXXXXXXXXXDDDDDDDD44444444GGGGGGGGGGGGGGGG4GGGgggEEEEAABBBBBB77766^^^^kkoo55aa0q�삉�~?O�r�3`�d�>���Ɏ	#���.�'�} }O�d�y�y�y�y���}DRPt|��N�/�G
1d̑�g4�/�(>#�'����05Hookk^^^^^66666777BBBBBBBBBBBAAAAAAAABAAAAEEEBBBBBBBB77777777BBBBBBBBBBBBAAEE77777777BBBBBBBB7BBAB767777777766666666777777777777777766666666666666667666^^^^^^^^^WWWWWWWWWWWWWWWWWWWWWWWWXXW9WX<DWWWWWWWWXXXXXXXXXXXXXXXXWWX<<XWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWXXXXXXXXXXXXXXXXDDDDDDDDggggggggggggggggggggggggGGGgggEEEEAABBBBBB777666^^^kkooo5aa0q���AD�F?����pY�i�>Ϸ����#���H��> <\ �� �X���>����}c�2x<� �@�"���;��S�G�1d̐=>٧�~A@���Q(�O���	�C{[Z�����������ٱ�������









***���������


)�����������������
��ٹ�������������������������������������������������������������������������������������������������������������������º�����b���������������������������������������º������������������������������ʺ��������������º�������������������""���:::***********************+;:***


���������������[[zA��	�����d��>
|AM�6f�����Gϓ�����Px�U�,�>a��E(2]��>�����O8�����p'f�#�ď�H�g�4�/�(>F?N%� ��0a5HHoookkk^^^^^^^^66666666777777777777777777777777777777777777777777777777777777777777777777777777666666666666666666666666666666666666666666666666^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^XXXXXXXXXXXXXXXXXXWWW999WWWWWWWWXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWXXXXXXXXXXXXXXXX<<<<<<<<<<<DD@@@@@@@@@@@@444GGGgEEEEEEEEAAAAAAAAEEEEEEEEEEEEAABBBB777666666^^^^^koHH55aa0q��C �Q#O��
nY�i�8H�HpJ	>DU����_�� �p	�Y.��'��	�φ|3�@��>i�L�"�:8p2*|�	>,�=Ji�n_��>D?N%����0aaHHHoookk^^^^^^^^666666667777777777777777777777776666666666666666666666666666666666666666666666666666666666666666^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^XXXXXXXXXXXXXXXXXXXXWWW9WWWWWWWWXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWXXXXXXXXXXXXXXXXXXXXXXXXDDDD@@@444444444444GGgggAAAAAAAAAAAAAAAAAAAAAAAAEEAAABBB777766^^^kkkooH55a00q8��AĢ~#O�rܿ-�-�8O���>G�\����*��4��~)��O�;'��8yߋ>��>d��O���I��3��8PY3�Je�n[��D#�%�Őq0���$7������������������������������������///////��������������������������������///////////////////////////////////////////////////,,,,,,,,,,,,,,,,,,,+��,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,+������������������������,,,,,,,,,,,,,,,,,,,,,,,""  #������������������������!!!!!!! �����������!���������/5����������8�G�A��Q?���Źn�fO��d�����8>��|�|�(<,��~���R���~�2��d�<��2v|2�5���d����8��#�Gً$d���p[��������q?��MMMR��������ח������������������������������������������������������������������������������ח������������������������������������������������������ח����������������������������������������������ח������������������QPPP���������������А������������͍�����ח�����������XXLG�� �q(�H�@�)�n��e	�c�G�p�(�O2q���~-��N�~<�,�Y~6�@y���|
���'�d��8�J�I@C��W�#�Ř�g�}�Lۂ�?/�|�F#��A���aaa555HHooooooookkkkkkkk^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^kkkkkkkkkkkkkkkk^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^kkkkkkkk^^^^<<<<<<<<<<<<<<<<@@DDD<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<XXXXXXXXXXXXXXXXXXXXXXXX<<<<<<<<<<<<<<<<DDDDDDDD@@@@@@@@444GGggggggggggggEEEAAAA7777777766666666777777777777666^^kkkkkkooHHHHH5aa0q8���A��Q?��@����6ͳ%z�C�Gϓ�	���2U��"���;>�����ә,���G���_���e��%��~��O�.|�O2T����م�H�A8,Œg-�p[�����Ő?�0�����$$$$$$$5��������///////////////////////5������������������������������������������������������������������������///////////////////////////////5��������///////////////////////5��������������������"""""""""""""""    """""""""""""""""""""""""""""""""",,,,,,,,,,,,,,,,,,,,,,,,""""""""        #��������������������!!�����///5��������$$�����8�G�C!�q(���b1>
~[���$[�|,�����"�p�~ y8���~�����Gc0;��_��,?�~2~���%������\�A��G�C��S�Gω�d�Y��ٶ�|AA�!�~(����������������ս�������������������������������������������������������������������������������������������������������yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy��������yyyyyyyyyyyyyyyyyyyyyyyy��������������������������������������aaaaaaaaaaaaaaaaaaaaaaa`�����������			����������������������������llmyyyy��������!! ���Մ���?��D�F#��@S�ܷ4}����3�G��\�����>���;d�� y����<�7��ǳ���,3f
�x�C�(������O2T�O����H��8,�=>٦i�p[���Ȅc�D��?��N#SSSSSSSV�����������������������������������������������������������������������������������������������������������������������������������������������������������������������涶�������������������sDC�CDCDttsDDDC���������DDDDDDDDDC����DtsDDDDDDDDCDDDDDDC��Ņ��������DEu�SF�s���������DDDCE�vtsDvtttvvtTTTTTTTTTTT$$$$$$$$$#sssq�����������������������ᱱ�������涶���􄄄�SV��?����D�~#�@���nm��!�$f'Ď>	p�| x� �G�'l���l< �Y,2X~9d��p��p})��%7����~6�����s�2y��RGG��/�G��1|%	�̳Lۂܿ/�(>#�'����000aaaaa555HH55555555ooooooooooooooooooooooooooooooooooooooooooooooooHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHooooooooooooooooooooooookkkkkkkk^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^kkkkkkkkkkkkgG@D@g7^4444GGGG444@@DDDDDDDDDDD@@@@@@@@@@DDDD<<@4GGGG4@DDDDDDDD@@@DDD<<DDD<<XXXXXX<<DDDWo@lDG<<<<<<<<<DD@@@4444gAEG@@4GGggEEEEEEEEEEEE77777777BBB77766^^^^^^^^^^^^^^^^^^^^^^^^^kkkoooHHHH55aaa00q8������q8�O�b1��-�p�l�4}�����8�'�DtE/�d�'.�Y�Nf~��M�����w_�O�o�G����_d�G}��%��~��@�8� Q@C��	(,��'2����~A@���Q8�O�'���������������������!!!!!!!!����������������������������������������!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!�������������������������������������������������������������������������������������������������������������������� �������a���aaa`���]m��� ����������������������lmyyyyyyyy����������������yyyyyyyy�����!! ���Յ�����q8���C �q(���b!��-�p�`�h�|,����E\� . >���'A�Y�+%6JDw_�L��-"�%��ك���~>�����%����	����> �	�H�A8,��8Nh���
Ȅc�D�?��N#SV�����������������������􄄄���������������������������������������������������������������������������������������������������������������������������������������������������������$$!��cEtTTTTVvvttsCCCCCCCCCCCCCCCCCCDCCCCDvvtsCDDDC��Ņ�DC��������DD�TEtD�CCCDttvtT$$TsFtTTT$$$$$$$$$#cccccccccca����涶��������������������������������􄄃SSSV��?���D�~#����~[���ْ��3�Gϑ��	�K%\|�O��d��!@����_�_$w�~ ~;?��#������o��,�Y��~���|��2T������#�Œ���̂ٶ�~_P|�F?J,�A��q8�N'����������������������!!!!!!!!��������!!!!!!!!!!!!!!!!!!!!!!! ��������������������������������!!!!!!!!���������������������������������������������������������������������������������������������y�!�l���		��� ����������������� ������������������ٽ		���������lllllllllmyyy���������������������������!!!!!!!!!!! �Յ��������q8����!��8����1>>/�r�8,�,p�l���<�'�G�}A�}b(�������������양�}s���v���v"�0!�����O�A�N(��@�N :>s�>Dx��`��8Y�i�n���|AA�1��Q8�Y����?��N'���
BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA��������������������������������BBBBBBBBBBBBBBBBBBBBBBBC{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{[[[[[[[[[[[Y��`�ll�¼66ln��������������������������΀�hh�Ί�h�Ί�Ύhhhhhhhhhhh������h������xx������h����h���hhhhhhhh����Ί���Ί��n�`����nnnn6666666666666666�������ސ�����������������������jjjjjjjj�jjj����```�q�������d2'��D��O����-Â͂٣�=d�Ġ���f> �d��.�Py�2P�`<��ҙ����#��iH�E(�Z}q_$wO��#�%��|6K�	��P �/�G
1|'��p�Lۂ�7/��
�����q8��� �?��N'������������������������BBBBBBBA����������������������������������������������������������������BBBBBBBBBBBBBBBBBBBBBBBC{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{[[[[[[[[[[[[;{ �քn��ּ6ln�������������������������΀�h�Ί����Ί�Ύ�hhhhhhhh��hhh���hh������������hh���hΎh�����������Ί�������������nnnll��������������������ސ����������jjjjjjjjjjjjjjjj��������jjj��````�q8���� �d2�ČF"����~_��f�l�4}������8E\���<Y<�?���e�f�{~
�
Gp�$Q"�H�E(�D�$Q#��w>�}|<`��s�\�N >��0�	#�Œ'�����~_�>D#���D�qd2�C �?��F����������������������������������������,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,&������������������������							��������������������������������������������������������mmmmmmmmmmmo���1E������xl����			�������� ��		���������ѝ������� �������ll��m!	������yyyyyyyyyyyyyyyy����! ��!!!!!!! ���������������Յ��������Յ�������q���C �d2�ČD"�O����-�r�`�i�>�1($|�Wp�O2p�L��~k�`��g�ߏ��}q���\Gi���\�iH�}<��%&`��J~<��d�� }O�>�|�G�$(O����-�r��/�(�F?�%�D�qd2,�C �?��N'���q8�MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXMMMMMMMMMMMMMMMMMMMMMMMMR�������������������������������������������������������������������ŝb-F�!ټ��j�ln�n�n�ւ�lnnn���������������������������Ύ�����������������Ύ��hhhhhhhhhhh��������Ί������������nllnll��޼�������6����������ސ�����jjj�������������������````````````````````````�q8�N'��?�����F#��P)�n[����L�2p��E\���N ��<���vN�?~�p��~9~
�
E������d���(�D��;H������`���������l�>��������|H�,�fAnpܿ/������B!��Q(�N'����d2������q8�N'	������������������������
BBBBBBBBBBBBBBBBBBBBBBBCzCY�Y��{Y����� ս�!!!�lٽ����������������� ��!���yy���y	����08\%��nqn�y���!�� m		x�����			�			�������������������				����	��y�yyyyyyyyyyy��������!! �����Յ�������������������������������������q8�N'��?��������d2'�D�F"���n[����L�2p�lď>	|�>s�>� X�Ň��6J�3~>�p�z#��k%���Z�k%���Z}q��Qf�t}y�#0�a�~�[%�8� �#��p"*|���>$Y}� ��n_�����B!��Q(�N'����d2������q8�N'��������	������������������������
BBBBBBBBBBBBBBBBBBBBBBBCY�@��Y�Z�Cy������zA�{{{{{{{{{{{{{{{{[ZA���Cy��j�ll������,JJ�^a?�$��!�S��cccst$$$#csst$$$$$$$$$$$$TTVvvvvvvvvvvvvvvvvtTVvttttttttttttttvvtTTTTTT$$$$$#ssssst$$#q�涶������涶�������SSSSSV���q8�N#���?����C �q8�J%1��Źn[��3,��E�bGϓ��W>�)d��O�|3��d���07��ҟ�ϧ��Gi�Q"�%���Z� }qY���>���#��Y?~,�L� �#��p*G
	�8$YB}� ��n_�����B!��Q(�N'����d2������q8�N'��������	������������������������
BBBBBBBBBBBBBBBBBBBBBBBB�Y�[z�BA��[ �!���!������������������my� ����!����� �����\ �u���^L��1E��ll�`�o7666777B66777777777777BBAAAEEEggggggggEEEEEEEEEEEggGGGggggggggggEEEAAAAAABB777BB777666^666^kooooooookkoooHHHHH555aaaaaa00q8�N'���q8�N'���q8�N'���q8�N'���q8�G����?���C!��d2�ĢQ?��b!>
|_�n[��3,�z������*�'�|R�W �1���P;�`o�Ϧ��O~ >���;H�EKY-~ >�����������������ed�y����	('��e	�̳nr��/��
��c���Q(�N'�Ő�d������q8�N#�������������������������@��Z��{	�BA�"L�͗������������������ך�XXMM���MMR����ဎ�G�+�IΈq�$GY�󈌼��666ll��666lllnnnnnnnn������������������������������Ύ�������������������nnnllnnnll666j�����ސ����������ސ�jjjjjj���`````�q8������q8�N#���?�������?�������?����C!��d2����q8�N'�D�~?��b!>
>/��ܷ-Âf��e�>��	88:�>�%ߊd�<��a���|�Q�������GiH�E(�\Gi�����W�`��J~<��d�� }G�|���$x��LP�g4ͷ���� ���F#���D�q8�N,�C �?�������?��N'���q0��������������������������������0������������������������$$$$$$$$$$$$$$$$$$$$$$$�����כ�L���`�6l������������������6�ސjjjj5kHq�F�` ���AX�(	#������-f��������涶��ᱱ�ccccccccst$$$TTTTTTTTTTVvvtTTTTTTTT$#sssssscca�cca�������BBA��BBBBBBBBBBA���	�����q8�G����?��������d2�C!��d2�C!��d2�C!��d2�C!�Q(�J%�D�~?��b1�D��O����-�r�8 �i�f_�|,���#�p�>�p����Xy��(���K�����-d���(�D��;H�"��`B;ρ���C�C��|��?�N����H��d̘�>�i�n�����B1�~?J%���q8�����?��������q8�N'��````````��������������������������������````````````````````````������������������������������������������������j�`�05HH5^7kd�7���0�7��������������������7��L��LR B@��b�88 p�q!J)��?0������$$7������//�����������! ���!!!!!!! ��������������������������!!����������///8�R��MMMMMMMRMXXXXXXLN'��?���C!��d2�A��q8�N'�!��d2�C!��d2�A��q8�N'�D�Q(�J%���F#��B |>>/��ܷ-�p��٦e�(J��<�$U�Ϝ��<�8��'o�C�d��<�����'���D��럀��~3~
}}�#0�Gӟ�vP#�x<J ��O�Af,��'�2p[������!�~?�%���q8�Y�A��d2�C!��q8�N'���q8�N'���aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000000000000000000000aaaaaaaaaaaaaaaaaaaaaaaaHHHHHHHHHHHHHHHHHHHHHHHHok^H(�'�V���cu����V����������������VT���&�f�W��������� �u��oqp�J���LXXMMM[�����ח�����������А��PP��������PPPPPPPPPPQQQY��PPPPPPPP������͍͍����׆��ח����R�����MMMMMMMMMMXXXLN'��?���AŐ�d2�C �Q(�J%�D�q8�N'���q8�N'���q8�N'���~?������F#��B |>��n[��pAl�2̳G	B�N	#�Ȋ�	�>��d���?|
}8���&K��ǌ���v`���->���������k%0�C�f1�+'l�d�yQ;��	�(,Œ2C��fAnr�� �P|>D#����D�Q8�N'�!��?���C!��d2'���q8�N'���q8�L,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,&,,,,,,,,,,,,,,,,,,,,,,,)																								����l���llj�aH5ooHHHk6oooooooooooooooo000aH^67F}�Y��#SSSS����Qqq`�����[�� �{�����h�jl��#����7������/5������������! ����������������!!!!!!! ��!!������//�//5�������$�������8�XLN'��?�����q8�J%���~?������~?������F#��b1�Q(�J%�D�F#��b1�F"���|�D"�B!
���~[��pY�X,}�!�$8%�Áp�(�#��G��ӈ�f������ǌ����v`��ك�?>��}�#�B;(d银O���J��;��R<pY zE�'2p[���"�b1�~?�%���q8�N'���qd2�C!��0q��#S���q8�N&���q8�N#���q8�N#SSSSSSST��������ST�����􄄄�����ScT�Q�T�����F��������q��������CzA�	�C�ռ��u�ܳ���RO��E��Ĥ���w�������?�`� ����s�6��8�MMM[ך�����������͍��͍����А�������������������������P�����͍����ח������������MMMXXXLN#��?���A��q8�N%�D�~?������~?������~?��b1�F#������~?��b1�F#�B |>
����|>��@���|_��n����g�B�FbPH�"�ptE. d�%ߊ;�B�ߍ?f�|�Y���w����f ~
��M������;�Ed�'��P �L��$}��,�8Y�h���D"�b1��~?J%���q8�N'����d2�C!��?����	�����������q8�N'	�����������q8�N'�����������q8�N'��������	��������BBBBBBBA��BC{{{{{{{{{{{x���y����`l`�q5����������$5�����7��$$������ۭ�{�qd8��%���Ĥ��������Ǣ�.��GҲ"AE�n'���Ž������!yyxll���ll������																										������llmyyy�y�������!! �Յ��������q8�N'��d2����Q(�J%���F#��b1�F#��b1�F#��B!�D"�b1�F#��B!�D"�@�|>
����|>��@�S���/��ܷÂ͂�`���"�1>$|�W>s�|��|�O��d��6J�~������씏�M>�}(����`���?~�;'g�>a���������O�Ad��P�,�4ͷ�����B1�~?���D�q8�N'���q8��C!��d��C ��000000000aaaaaaaa00000000aaaaaaaa0000000000000000000000000000000000000000aaaaaaaa55555555oooooooo55HHooookkkkkkkk6BHq$����R�+��������m�&��&A���05k0oa8��U�B���"�R�F�(hf%秥�ǧ���Ĥ��������[����	��7 �!E�jj`HHHoooookk^^^66777BBBBBBBBBBBBBBBB77777777777666^^^kkkkoooHHH555aaa0000q8�G����?�����q(�O�����~#��B!>�����|>�����|>�����|�D"�B!>�����|>��O�����@�P(
���~_���n[���f�`�Y�p�/���G߄�\������DP�/�߃d���0;���)�Sd��}��0V`/Ɵ�����C�\�A��G����������fY�[��?/�(�D"��c���~(�J'���q8�N'�Ő�d2�C!��8�N,�����������������������������������������������������������������������������������������ս���������!!����yyyyyyyy�m�!���ݬ�x��m myyyyyyyyy�!�xmy��q0���$8�����Ȍ'�A��~d�A����K�OOOOK��II@ E�E����/��p8����>'��ST�������������ᱱ�cccsssssssssssssssssssssssssccca���ᱵ�涶�����SSSV���?���C!�q8�J%���~?��B!�D"���P(
�@�P(
�@�P(
�@�P(
�@�P(
�@�P(
|_��~_��|_��|_��~_��n[��pY�X,̜'�z�	�('Ȋ��@?���(�A�|�@�v?�#00�C���`$va@��~)���d������_��L�'���ٷ�|A@�!�F#������Q(�N'���q8�N'C!��d2�C �q8�N#SSSSSSSV��������ST���������������e�sfQ��T��v����������d#sf��ce�S�D�~#���7�ca�>j��H��EEC#$3��������P�aq`�c�0������s�A��?$B���`�jj�������ּ���666lllnnnnnnnnnnnnnnnnlllllllll666�����������ސ��jjj����``�q8�G�����dN'�D�Q?��b1�D"����|>
>/����/����/����/����/����/����/����/����/����/����/����/����-����/����/����/��ܷ-�r�76�٦d�"�18'Ď>0���2T�G��O��t��s%���~0 x��?d�c�G���~)�����RP �o�G��d�Y�p� �m�n��>"�b1�~?�%���q8�N'���qd2�C!��?��A��`````````������������������������````````��������````````������������������������jjjjjjjj��������jj�������������֐�n��^68��LO������������f�#��>Q8��L��D�ѐ}���2P �����`deEC$3����c"��qqaaqaaqp���x����
?�'A���HHoookkk^^^66777777777777777766666666^^kkk^^^kkoooHH55aaaa000q8�G�����dN'�D�~?��b1�D"��P|
>/����/����/����/����/����/����/����-�rܷ-�rܿ/����/����/����-�rܿ/����/����/����-�r�7-�p�`�X,�%�d�����8ap�| x�����P �w��?c%��A������;�/Ŕ���#�(�>s�~>|Y�zP�,�2f���ȄB!�F#����D�Q8�N'���q8�N,�C!��d2#���q0�0������������������������0��������0������������������������������������������$7�����������������Y׏�fē�B+[[[[[[[[[{Y�:"��F"�'����KzȲc�,��-�
V�(�#*!���!������������=�@����X����
����!!!�����yyxlll��������������������������lmyy����yy��������Յ��������q���C!�q8�J%���~#��B!>��@�P(��/����/����/����/����/����-�rܷ-�rܷ-�rܷ-�rܷ-�rܷ-�rܾ/����-�r�?/����/����/����-�p�7-�p�`�X,�%�d�����EY��Ϝ��<C��G�"�'��H��'E?k�o�
(���_�>@��}g �T�H����"�pY0z}�,�2ͳm�r����B!�F#������Q(�N'���q8�N'C!��d2����0a500000000aaaaaaaaaaaaaaaaaaaaaaaa00000000aaaaaaaa00000000aaaaaaaa55555555aaaaaaaa55555555aaaaaaaa55HHooooHHHHHHHHH5k0q/�9�ȇ1B+{{{{{{{yD��4��ҀjD|C�`���c�EJ0�e���7�rddddddddeEEEEEEED44444442���qg��1��u�   � 2���l�� ����Մl�y��ݝ�լ���lmyyy�llllllllmyyy�������! ���! Մ����0q8�색ĢQ(����1�F#���|>
���~_���~_��n��n[��n[��p\�p\�pY�m�~AL�
n�i�n[��n��n��n��n��n��n��n[��n[��n�pAl�2}����3�PH��"��G���d��Y8|�K�\�oŲv�	��H��,��K�q�!�E/�>�p2*�$p��LE�,�,�������B!�F?������~(�N'���qd2�C!�?��N#���q8�F,,,,,,,&��������,,,,,,,,,,,,,,,&��������,,,,,,,,,,,,,,,&���,&	���,,&&�E�y��l�58��J&�f�g�����#��#P�DiDX�̡?�W����� ��l��M���y��qcV��TQlQ� ʉ�(� z.db��(������������������y�p��s�$$$001� � 9^5dY&deᴃ���� �	��lllmyyxlllllllmyyy�������! ������Մ���?��G�A��Q(����1�D"���|
>/����/��ܿ-�rܷ�p��p�7�p�3l�6ͳl�6͸,�4̳@��>ۇ��f���p\�p\�p\�p\�n��n��n[��n[��n[��p\��L��E�HɎ	�#���Y��\����*���2p���('��>�φ|0�|P"(2q�̕���80�	�#��B,�f�`��n_��>"�b1��~?����D�q8�N'�!��?������q�����``````````��������jjjjjjjjjjjjjjjj��������jjjjjjjj��������jjjjjjjjjjjjjj�jjj���`l�qq5���M������4aEx�[���G"*̤��D�����oB{*����1#�D�x\�dؾ,��s4>��C1*�<R�**����*������������������������d��^z\J.,�{��Ꮀ��!a';b;y��j�ld��!�f�涱�csa����������������涶����􄄃SVV���?��D�~#��B |>�@���|_���~[��n��n�fٶm�fٶm�fٰX,��`�i�8O���f��m�pY�e�n�m�fٶm�fٷ�p\�p\�p\�p\�n��n��n�fٰ[4̟ez�Y#18%�?	fp#�#�)~#�ɓ�>�'�|��0���d��� �|�;��S�G���dτ�fA`�m�n��"�B1�~?������Q8�J'�Ő�d��A��q8������```````````jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj��������jjjjjjjjjjjjjjjj�jjj���ސjjj���`�j��j�?������eW�{�>�����/���"��T���� �:@i]���\�$ͲGJTd�@�BL_� gE%\�*c�خ*T�D
�TTTTTTTTTTTTTTTTCCCCCCCCTT2C1//=...%%%{�ÉE�o10'���䬈�`�`FH^6ka0o7^^^^^^^^^^^^^kkoooHHH555aaa00000q�����Q(���B |>��@���~_��n[��n��fٶm�fٰX,�3@�X,��l�4�3L�4�3L��p�g��}� �Y�� �Y��3L�4�3L�4��`�X,ͳl�6ͳl�6�7�p�7�p�7��l�6f����"����3�G���	p78:"��~#�*� �p�\� �y����S�(�8p"�ȏ�ə!p�@�m�n���Ȅb!�F?������~(�N'���qd2�C!�?��N#����0000aaaaaaaa55555555HHHHHHHHHHHHHHHHHHHHHHHHooooooooHHHHHHHHHHHHHHHHa55HookkH555aaa0q8�A�2����QHzn��m���{���@ Ou	=��˔S'1{�7����IKTPm2,^�pt���O�a�銐&LQ���)*RJ�Rdddddddd������������������dd��bbbb^^zzzz^\,�./O2=.=111`/s�$���.&�a��������ᶶ����������SSSV��?�%�D�~#��P(��/����-�p�7��l�6͂�l�4�3L�4̳,��p�'	�p�'	�p�'	�p�'	�p�,�2p�'�BP�,��� �YB̳,�2̳,�2�3L�4�3L�4��`�X,�.��.��.�ͳl�,�3L��}�$[$d�����<|�����A> �H��O����p� �W�?�����>wf�|�G�	�f/�=>ِ[6ͳm�r�� �!�D"������~?�����Q8�N,�C ��d2������q8�XXXXXXXXXMMMMMMMMR����������������������������������������MR���MMXXXL�@��!ĈDy�7����'�Dࢅ|��?֨� 

���B�;1Akq�}	�Z��(��T��'��O\TPq,�ҡH` �)2d	�Rt�U)����������������̌�����LP�LLK������������w��X��Y��../. )<d�K�T������������􄄃SSV���?���D�~#����)�|_���n[��nm�f�`�X-�f��e�8N��8N��>���>ϳ��>ϳ��>ϳ��>ϳ��8N��(C���Nh�8Y�Y�}�g��}�g��̳,�2̳,�2�3L�4�3L�4ͳl�6ͳl�6�.6͂�`�[4�3'	�}�o��FbpJ	#ςE\�� ���� }G�}G�}DRE/�(�8p7�~8Gϋ1d̐�(Ni�p\�~_�P|�F#�b1��~?����D�q8�N'�!��?������q8�F,,,,,,,,,,)															mmmmmmmk��������mmmmmmmk��������mmmmmmmm��	���)���,,&	���RAEx��E/O onY#��@�QT����V�%
��4��(���d
�)\��t�4�"eJ�2CLuIԬW&t�өT�\�*�Ɍ����������������LLLLLK���LLK���L���Q���K��̐��A����E�^oH,&��'�	�C{zBBBBBBBBBA��	������?����Ģ~#��@�)�|_��n[��n�L�4̳,��p�'��}�g��P�%	E�dYE�dYE�dYE�dYE�a�P�$[�f'����"��(J��(J��8N��8N��fY�e�fY�e���`�X,p\m�f�`�X-�f��e�8N�=|,����PH��|�p7pp#�>��#�:#�:>�>��>w8*G�>,œ>�P�,�-�p\�~_P|�F?�b1��~?����D�q8�N'�!��?������q8�XXMMMMMMMMMR�����������������������ח����������������������ך��X\G��A���	���Y$،����^Ӏ�_O4V���T��9P�S��ɣ'�\bb�۲b�H&
�إ�X	����R	�*�s)��Ru*eɓ1J�2c#######%EEEEEEED44444442�������������B�qar�Qs�QqrRQp����p��I�{ͨ� ِq0��7�$$$$$$$������8�N#����8�J'�1���O��ܷ-�p�7��l�4�3L�2p�'	�}�g�BP�%	BP�dXz���z���z��YE�dYE�l������f%�Id����bpH�,�"Ȳ,�"���8N��8N��8N��8A`�X,��m�f�`�X,f��i�fY�,=|,��3�pO�A#���$T��Vap7>s�8�>wp'p8�>D|���ə#�O���f���p_���Ȅc��F#������~?J'�D�q8���!��?���'����	����������BBBBBBBC{{{{{{{{[[[[[[[X������������������������[[[[[[[X��y����QH555aaa0}������6�r�2 %P2
*{P�r�ǥ���\�b�)rU�I�uHWjB�!��b�Y9jyR��� �)�J�Rt�d�S&..==/1CC=12TT21=/1C2TTTTT2C1=.%%.=1CTT1111111111/=%==.%%{��:���C���A���jּ~68�������~8��G�AD�F#������-�rܷ,�4̜'��}�l��}�,�,�"�3$|!�z��P�l���b��>ɟ	Bp���fbpN	�8'���H�O�$q 7�ٳ��ql���">Ɋ�=C��(O���(C�,�>ϲ��8Ne�f�`�i�f�`�m�f�`�X-�fO��="���|,���>G��>G��R*EH���	����	��	�#�x����Y zP�g4�np�7�����@��|�D"������~?J%���qd2������?���'���q0���������$5���������� ������[����͍���א��P��������Й͍�RH(&��cA���A�ݬՄ���
sFP4q0�#��,",A�RaB�*T�RX�*L����T�J��ӪT�:T�2eN�:�*U)R�J�*T�H)bu0�X�:������ȼ��QP�ļ��X88��Qļ�������������������ļ���\\�����\\X\\\X9��G(����EĐ���(�W�L�C�D���Մ���O���3`��n���϶e�n�m�8Y#�H�,=|/��"Ȱ��c�|O��>Dp��bɊ%-�H�$8'���b�a�&f,��"MޞN��%��� ��#�rp�B�G�&J�=d�Ċ�`[6P�`��>ϳ��fY�h�3L�4�l�4�٦d�>���"����Y!�>%���<G����	"�T��	�#�|���pY3$J���ٶm�n���|_P(>��b1�~?���D�q8�Y�A��q2������0q8�XXXXXMMMR��������כ�ך�ЌF��RF͍����Й�M�ח����QR����#dsSd��R��A�q(�/�ؘ� ]��q9"�$.R�@8D�z��b�*L�Rb��L�3�X�ӎ�R�*S�N�J��Ҥɕ:t�T�T�J�*T�R�&��U��):UI������y����y��c��\dzz^^^bbbzz\JJ.,,zzzzzzzz��b^z\\Jz\\\JJ...JJ.,�	QPeg0�&�mm��l$c�CyD��~(�N%0}�~_��
|_��|[�Y�E����E��G��H��d̘���>pY�m�8H�H|J	�8��U@���4DfH��8J(G+���Fjp'I����}�<��I�J�#9�"�	f'�6}�B�PY!�̳$YBP�g2̳L�2̳L�,f��X-�fN�8H���_zE�fL�N	�>%���>G��#�p�"8G��A>'��L�҄�8Y�[6͸-�pܷ/��
�����F#������Q(�N'�!��?���'��q8�XMMMMMMR����������כ�N&�sv�sctT�ccsst$$$d$#d$$CE�$���!���6`�7Go#?'��Fl��� ~��^W{�%*��9H�eE':LP�d�&L��ʝ&t����)R�:t�T�R�:T�R�N�J�*��R�J�*U$Ա:��bd222TTTTT1CCCCCC11% .C%=/11111////=........CC11//==......%%%%%%{�����pK�@��Fn[�ĈD0�����c��D��@�0}�n�n#$|!�E�%6}����CY����)�* h�t�A��t�@��\-K�� o������n�	�ĉo ��17؈�M��{�J>|����J	Ad�Xz���(J��8N��fY�i�f��e��٦d�f٢��@��8C���FLə�18'���|J	A('���bə#$|/�="ϳ��f��m�n���~A@�P(>"�b1��~(�J%�D�qd2�����q8�N'���	���BBBBBC{{{Z���������z�AD��l�n�����6nn�������n�h������ސh��lؐnn���~am^op����bM�/�c&��3�PY���$��`` T�Rb�&)8�ɕ:��RaS��J�)ӧJ�:t�ӧN�*t�ԩR�J�*T�R�*��X�``UQQQQ��ļ�\\�����%.=/%.=/1C22........1111////......==%....	==VDAgAq7%�}�8�O��,�0|>D#?,���_	Bn�QE!�U�U]�a���p����D�Og����}��B o!�S��$&�}��^�&�Ù��}:��bbo�Ј���{=�.�'ИC*C4PY���,�$#�x��G��C�,�(J��8Ne�fY���f�`�i�f[�Y��,�fJ��"����Y#�|,��2fLə3&d̑�>�=H���>�e�f��n���|A@��|>D"�c���Q(�J%����d2������q0��������$$7�7�������///////5���Z����ƨHCf���HHH((&��f�(�hH���$f�C�[��jx��`%mh?�����h(���(�000(�*'�'�QFT�Rd	�&��(Q�N�JT�1AB�*�)ӥJ�*T�ӧN�:T�өR�R�*T�R�J)4�GB��*�������dd�b^^b�db�d�d�^z�%.=/{�Åˋ�LK����������������K���OK�ˋ�OOK�Eß�/qs���D���ʻ��lnF~\D`�rͳ'2̳,�4���\��A�.�g؈���LLD	��p�����_o�����t�C@�����!�`�K� hi�"$H�t	��\/g���I��p��D�_ba�%�E�4�q>ȫ�����
&d̑�>�"ϳ��>���fO���f�`�i�pAl��P�g2p�'�BP�a�zE�dXz���C��="Ȳ,�(O���fY�hn��~_�
���B!�~?���D�Q8�N,�C �?��N#SSSSST����������������������&��V��e��[���������			��y]ax�����`�lD"6"��>�h�ޜ������J�d��=8�eF�D���&@�R	ʉ�
�:t�Rd&L�ӧJ�*L�R�N�J�)S�N�J�JT�R�J�*z{2q��N���#*!�����*�������������������������������������������ˋ��]d�������p�@�uy�pO�[�~?�8���\� �a�����|�CDD�O�����������{:�Ba�  �0ЇK��H$�}>���7S�E��}�8C^�g��i��t�>@�.���K��E��G�|Y�1f,��>��%	�}�g	�p�g�2��`�i��٦d�8Ne�8O���"ȳ�(J,�"�҄�(J��(Je�f��X-�fۆ�~_�
���B!�F?���D�q8�N,�C �?��N'���	��BBBBBC{{{[[[[Z������������ٳX�A����n�n7^B666777BkeY@ln�$>\�@NL��`����ؚ3�212d�$̓��`J���钡��ӓ§� (P��d	�*A=E8Q3�J�*L�2�J�:t�R�ɓ&L�өR�*t�ԩR�J�*T�R�OCQ`TO ��M*�eEC$45C#��%C����RT43###%ED43������������RRR�����RR�������������p����,�������M�/��Ѩh445��u		�]/g�����$$�}>�D��a7��M��{	�������`7�M�4�~�D��n'��DL45�&&�}	���_O�0�  �0�K���n�B��.�Ku���_ |���bə3$|/��(J��>���>ٖh��`�m��G	B̳'	�}�$Y}�g�BP�dYP�%	BP�%	B�3@�X-�fٶ�n_��
����!�F#���D�q8�N'C!�?��N'����	��BBBBBC{{{[[[[Z���������������X�Z�����;�ݬ�xlll���������q�Y��e`� uJ�t�q2T��eD�B���<�I�r20R	��	�***$U�
�(�eJ�Q1TO
L�Ҥʐ L�S�Ν*T�2dɓ*T�U*J�:u*T�R�J�*T�S̓£'N
U2��dddeC#$3���$3��3#���RR�5EC##$443�����qrRR����������3$c#�������RQq`��aa`���������  /�P� h�4&�}��o�����}��DDDDDDDDDDDDDDD^�g����{=���C\.��&"�}	:�O���DDDDDDDLLM��p�<�N�K���s+������$x���G���Y1�8,��f\h�"�e�|Al�4�3,��p�,�2̳,�2̳,�2̳,�2̳'	�P�'��̳l�6�.p�>/�����A��|>D"�b1�~?�%�!��?��N'���ս��555HHoookkkkkkkkH7ak76o56Ba<k7H?�4	A^o~Oȭ�!�d��Ѥ5�d�Y%1TF21=TFFFQQQQQON```NN
���(�E&L� ��� �)2��*L�T�c& �	�:u*T�R�J�)ӧJ�*L�ӧN�:u*�)��:T�U)�% ����(P���*u===EEEQP��ļ�����������������������ļ������������������������������\XX88XXXXX8889��{�����[�E�4�{	������DDDDD���a����{=��g�hhk��&"�}		>�o�1117����p�\/'����Ps:@��Pۇ�>w�d��$(Y1�f%2P�Fh�ٓ��٦i�fY�e�fY�e�fY�e�fY�e�fY�e�fN��8Y�i�fٷ�n���|_�
����!�F#��c���Q(�Y�����q8�XMRN&�ST���������������f�T����q�#DT#vT����L،jlʐ�H�h�u8ܖ_"B�䤈j��S�U��TS����Ә�
��+ R� L�AB�98)2X�*LQR��
NQT
QeN�J�*T�R�J��ҥJ�:t�ӧN�J�2e)N�&uJd�I�
(�B�:t�T������eEC$3���43������qr��$44444443�������RQqab���p��p�q�y��)(�����p���������pps����?��� N׳���}��������������������������g����{	����`0007��LE��}>�b""bbbbbog��5��p�:]#CCA��u��n�[�e.`�H�5�҂�?�S��'ȏ3�E�HpY��"ϳ��>�`�X,�3L�,��`�[4�3L�4�3L�,�3,�4�lۂ�-�p�>/�����A��|>D"�b1��~?J'� �?��N'�	�	�BBC{{{{[[[[[[[Y�zB�[z��Z�;yE��6�j\�  �ܛ<�_�b�7�1`��@�I���E
`QFOOONNN``N`
(��AE``
(�2dɓ&(+ QD�'
&@S �eI�*T�2S��
 L�S�R�J�*T�R�:t�R�R�J�*T�T�L�2��J�R�2R� L�R�R�R���999===QP���\��QPĸ\����XX�������ļ��ļ��\X88 $8����� 1�,\\\\JJJJ....,,,,....,,,�{����E�Da�og�k�	��}��Og����{=��g����{=��g����{=��""bbog����{=��g�hhhh���t�B/��u��s9��g3�i��PVP)s<���I���0��H�Y3&(Y�b�Y�&Nm�f��h��l�6ͳl�6ͳl�4�3L�4�3N6f��[6�.���rܾ/�����A��|>D"�b1��~(�N'���q8�F	��$���BBC{{{[[[[[[[[[Xۉ!�x�ٽy!y��A�B$C3d8����ׇ�4�"�/:,,��db�@��zrrz1��rs P�B�
@�2d

(QD	�:t�1L	��(�1AE*L�2�J� ��2eJ�:uJ�*T�R�*T�N�*U*T�R�J�Jd˓)Ju*�ɓ%:T�S�N�J�2d˘������TQ�����P��E�K��C��ĥ��&(hfFHhhhf&%��&%礢��� �bQp��  c�8XXX\\\\\���888XX\\�XXX889��������p�C���t��� oa0000000000000007����{=��a117����{=��bbbbog��4445��t�].��������s9��b�����������s����K��h5Y =>$p�\�_��_="Ȳ��8Y�e�fY�hfٶm�fٶm�fٰX,��`��f�`�m�p\�n��n_��|A@��|>"�b1�Q(�N'� �q8�F�$���	�!!��������������x����j�Gkg5?�����mM��;���|.I�swr1yz�%ED3%�d��eD46 �B�(P�eJ�&LP��B�&T�ӥI�`N L� �H&((��J�&L�ӥI�*T�ӧN�R�J�*T�R�*T�N�R�J�*T�R�r��R�L�2d�R�J�*�*S&\�r���������eEC##��5ED2�����W��8\�������������ļ����88XY� �u�:�@_�������Å���Ń����w��\Y���:�^O'����p�\.���{=��g���"""&&�{=����������g��45��p�<�CCA�����s9��r��33333335e�3u��s�U���6Tr3$d�(�~*|�&|!��d���p�,�,ͳl�6ͳl�6ͳl�6ͳl�6ͷ6�np��pܷ-����/��
�����D#���D�q8�'��```�Hoq3�8�������ך���������F׏�&���r��R�Qs����=�ٖ�A�!q�� �&I��F&I���aX������
(P�B��*T�2�@�R�N�*@PReJ�(�Rd*t�2ʥJ�)ԩR�:t��*T�R�J�*T�J���ɓ&L�2dɗ.\�JU˓&R�J�*T�L�r�˗.OOOQQQFFOOOQFTT2CCCCCCCC=/={��Ë��K�P̕�����LLLLLLLLLLLK˅��.�g����  u����������w�������=�BB@_�   !!��@3���y8\.���p�����������g����{	�����`07�hhk���y:]!����n���r��335eeeeeeeg%e���g;�ͩ���s/��Z�g�$($x��g�E�'��̳@�X,��`�[6ͳl�6ͳlۂ�`�[6�-�p�7-�r��/���� �P|>��B1�Q(�N'C!��q8�XR)������mmk��mmmmmmmml+��R��ˉ�>��`i2���>����b����)��F*�ʆH�����
QlB�((�ʓ&@�B�&T�2�J�&@�S��
*��D
�*L�3�T�R�J��R�:u2dɓ&L�J�*R�:u2dɓ&L�2��W&R�kɔ�L�J�)�.\�2e˓�TTQ�������Q�����̕�K�E��/������#%C##$443�43###��qaaas���3���y����������p�������@@B@_������=��`n        �������׳���{=��a17����p�@����CC\ @O'����t�_/��u��s������(++++++++9+++9=<59<5=��ܞ���C�Ҳ�E�#�Ɏ�"ϳ��f�`�X,��n��.��.6��lۂ�7�rܷ/����/��
�����D#�����qd2'������Ԣ���r������ּ����������j`�~"+ 	���� ��'�* �0��22 t����q1L	���(�I�X���*����(QAE&L�
(�R��*t�R�N�*@�T�H
 u)�d	�R�2d�T�R�)ө�&L�2dɔ�R�*S��.\�r�ɗ.b�2��X�L�2��T�L�2�ɓ&\�������������������������b,Jz\,��ŋѓ���Q����LK�K��OOOOOOOOE�������� q�	:�n��c�� , �u������!�� !� !!��!������X#�A�4�t�����������g����$�{=����CCCC\.���y<�O'����s9��r������5g''����������ׅg���5W�g����;�ɚ��ә����88EO�B�Y36̳��N	B�l���l�4�Gpp_�Źfٷ�����D�,���7$G�ܳ-�D�(����D�D~Yg� �D6555q��f�g��#x3K��6jjjQ?��7
��Ҡ��#���{�����(��!��*##(��#(��
 M9���(P���(� @P��H @�2eJ�*T�R�N�:t�ӧR�J�*T�R�J�*T�T�R�2d˓&L�2dɓ&L�2dɗ.\�r�˗.\�r�˓.\��+W.\�r�˗.bŊիX�b�999===EEQQQQQQQQ9ĸ����\X88\��D�QP���ļ�����������\\9��{�=�_�7�����q����  A�����:�a/��K� �� q���`a���444��{=��D^�`00���������y<�O'���444�|�\�w;�������AAY����ᩩ����ɥ����e��}��Uɱ�Y��饥AY̠�i4G2B<pH�LɊ�n[�l�,��8Ne�(N�8Y���fߗ�ܳ`�[����M�(>����B!��
���G�����R�s����^(��'�
�B;2� x}������a&Q0�tas�w�q)���y����2���2���2�{ QD�((�B� L�
�ɓ*T�ӧN�:t�ӧN�:u*T�R�J�*T�R�J�J�)�&\�2dɓ&L�2dɓ&L�r�˗.\�r�˗.\�r�˘�Z�r�˗.\�r�,X�Z��,S�������Q����������̋ˏK�K���OP�̕��Ǩ���K�OOOOOOOOOK�E������E��.��������u��o�A'Ӭ  %��   8�o�bA!00  '�44DM��p�\.���|�_-��u��s���%&ffj

�OOO----���-+,��+-��M
�-��-��L����MFfmג#rE_���R>����H|Y36��ْ��fJ��n
m�>϶�8_m�|[�i�?7 �h
���(��� ��(��~[�1��m5��-�&C����א�M��W�PawX��3�]P��J zdd���d��b^^�������dd����������S P�E
(Q	�&L��
 @�2eJ�:t�ӧN�J�*T�R�J�*T�R�J�*T�R�R�Jd˗.L�2dɓ&\�r�˗.\�r�˗.\�r�˗.\�s,V�\�r�˗.\ŋ�V��jլ	�����ꊊ���������������TK�ˌP�OK��LP��̌������LK�OK��OOOOOOOOK�EŅ��E�Ń�������  �	 y�:��`�� ��p�[�� �u����7�8����p�<�.������t��� @@O'����y:].�����u��n�[��3���s���������((99=<554������44/��������442�$���#������"/�2����J%��>٦bG
	�f٣�G�	#���F��!��=f��D���/�pq8AeP|��� �S��.	�|H�g��#��\�w%��fŕV���K�1�J�bJ\,J^� \z \z^b���bbb^^������dd�����������+ P�E
(Q	�&L�2
@�2eJ�*t�ӧN�:�*T�R�J�J�*T�R�J�*T�R�2d˗.\�2dɓ&L�r�˗.\ŋ,X�bŋ,X�b�s,V�Zŋ,X�bŋ�V�:իV�00''''��****************'0(�����!���������!������������������������������������X `K� � �t:b ��0w��� u�:� o��8����$�{8^CA��u��t�]#CA����n���w;���s�����((+((+++999<<54�����/��������*��,"��"�,""$��6  ��/6"���Z��Z�M�'$IH?���B3��Y���(Y��>ۇŹn_Ÿn\@��!�(�)pQnY��f��6��h�fJ��R��t8\/��3�08������9��=T.FT%F2%=111=.C112QOF2TTTFQOONOONN``
(P��
 @�	�&T�2d� @�2eJ�:u*T�R�J�*T�R�J�J�*T�R�J�*T�R�2d˗.b�r�˗.\�r�˗.\��,X�bŋ,X�bŋ+V�v,X�bŋ,V�q�Z�jЬ	���ʊ���������������H��&E���hhfFHhhhfJ��Hf%�秥Ģ��秧�������Ģ���� /��arRQarQg��9�����  /7�����bN�  �@   A��~�O�;���&�n���g3u��n�[�g3���s���%%&ffffffffj���NNOOOOOOMM--�+-�쪪��)))'�*�*�����(���i'#fȭn!����dC��0�kÓS��Ҡ���n���OMN,�>A���3$Y��8-��p�٣������8%�|[ג�� `��ܹ��u�:̋�BK��E�E�U�Þ�䤤������J�g�He�(fJ�HhfHfH�����*)��B�((QB� @�ɕ*T�R�ɐ @�2�J�:u*T�R�J�J�*T�R�J�*T�R�J�*T�R�2e˗1b�r�˗.\��,X�bŋ,X�bŋ,X�bŋ�V�8�X�bŋ+V�qݻq�
���998��������QQQQQQQQQ=99��QQQP��QP��ļ��������������\XXXX\\X9�,.J�{����w��� �8Ą�N�#���~���n78��HHH�~�] Ρ'����s9�JJJJJL����������������������ZZ[[[[VVZ�YURRR[NP�RV�Y��͐�ƕ��^��D��-�/�w���$.�X}����=��aM�,�
�(��1f������[����
(�1af%�jpPB�M�1 �����	%	��ÉK�E�	P�K����&E�ǥ��fG��&%�����*)�ʊ�,S�S�Ә�(P�B� @(QB� @�dɕ*T�R�ɓ @�R�N�:�*T�R�J�J�*T�R�2dɓ&L�2dɓ&L�2�˘�b�r�˗.\��,X�b�jիV�Z�jիV�Z���Gq֭Z�jիV�Z8�ݻq�
+rrq����������������z2�ql
��&J��(�ʈ��(ʆHhʊ�Hf&%秧������Ģ������e��w���c�9���Ş�w�c� %� ����`�BN�GC���t�>�N����}��O�А�#���|��9�((++++++99====99999999=<<<5554�������4,�4/�����666����+���3����!2�=<"?߭$�Ρ%�'�H���%�H�y�^bfa ��71{��"l_s*�9�K�Fe*|V����^BWt�?,��{P���Y�  �y���o��@ ���׺1y�������"���%E3 �	�*(ʈ�)��(���E0'�00@�dɐ @� ��
 @�2ɓ*T�R�J�&L��J�:u*U*T�R�J�*T�R�J�ɓ&L�2dɓ&L�2e˗.b�j�,X�bŋ,X�bŋ�V�Z�jիV�Z�j�+V�qݭZ�jիV�Z8�v�q��0��*)����F%��P̑�TTTQ�P�B���b����b^zbbbbb�dd^b����^^dbzJJJz^\.,,JJ,�%..	{���`   /���889��		:�_�/�@S���t:D�߯��P83�4I��$u>�_BO�ۨ���zxhejxjrs�=95554==<<<5554(=,�<46��94������*��,���#��7�:\O@� mOCO'���$�u���:�`/w��$1��u��b�C���u	��>��O���E��$u,�`��CRؘ8�3�!��q�����n0@@ [���	{��ÅˏK��LK��K�P̌������������������ӓ��
(P�B� @� @�
�*T�R�J�*T�R�J�*T�R�N�:�*U*T�R�J�*S&L�2dɓ&L�2dɓ)J�*U)�.\�r�˘�bŋ,V�Z�jիGq�q֭Z�jիGq�q֭Z�jի]�v�۷n�qΓ����������zd)=��<��E�(P�fJ��Hf%��g���*��(fJ�ʊ�E礢�ħ��e����礤�Ǧ/����$1��	���?��w�H```HH H  K��A��~�ā��C� �HI��q��O��k��&�t�Օ��Z�[Zڞ�[[[[VZY[W�RYUVRYZ�YZ[Q��^��-��gA�tYDI��q�:��.�p ���X#�%��	u��n�X  ���  �t:���o�b@a!'�����_ju���΁�� �  u�� @_�w�p��p�)�y�����y�������������������zzrrs �B�
(Q @� @�R�J�*T�ӧN�:t�ӧN�:t�ӧR�J�J�*T�R�Jdɓ&L�2dɓ&L�2d�R�R�3,X�bŋ,X�bŊիV�Z�h�8�:իV�Z�h�8�:իV�Z�k�nݻv���:���0
�(Tc�6i����ʌ���)��#(����*'������TFQNN`NN1/..=12F21=/11/.CT		{�?Ï_��F!��!�����/�X�K���~�:����N����t?IC��7Q ������}���O�7И�Y��U}AY�]��%}�ee}U���U��U�������}�\�	a��3 gy�
2{�ˏCC��3�ac��续� ���:�n����8883��$$H�t:	N�w����q���ď�G�%�� y��?�CBB@@@C���������OLP̌����̕�TTTTTTTTS�������ӓ����(P�B�
 @�&L�2dɓ*T�R�J�:t�ӧN�:t�ӧN�:u*T�T�R�J�*T�L�2dɓ&\�r�˗.\�JT�S.bŋ,X�Z�jիV�Z�jիV�q�q�Z�jիV�q�q�Z�jիV�v�۷nݻq�\�� ��*L�T�%iE*���NQFQ` u��(P�	�)��f&*��	��H&L���22� �he�ǥ�'��Ī,���/��[���.C`Q	��?ş� ����gP`�@@���	t?TK�@���"@�"O�'C���}>�Bo�5�ˡ���Ъ��ʾоʪ������������xrx���r��r6ֲ�$Q|��=�L�ş��& ����a$��'��.�XHs�$0000$0��~��C����$t:����"G��I��t:��N�����u:���@w���u��À@_������..%%.=12TFTTQFTTTQONNNNNNNNNNNNNNNNNN```
(� @�dɓ&L�2�J�*T�S�N�:t�ӧN�:t�ӧN�:t�өR�R�Jdɓ&L�2dɓ&L�2e˗.\�r�ɔ�R�2�,X�bŋ�V�Z�j��q�q�q�u�V�Z�j��q�q�q�wnݻv�۱�u��� L�RdΥ&�M�����������ɕ&@PU�� �	��	�:�*T�B�0&�J�����1���#���H���	F&(�8X��X�zd^,Jd�\.�u�8�o�� IU@g(�`8�����3�I�"�q�	8�^�/"B�璃�CbJJJJJJ��*�@��9�:�b���cu���ҲH�`O	.FOQ2.����E�����K�����q`�HK���~� �7@3���t:� ��Q ;��I�H$"�q� 8�`��[���%//==..%%=/CTFQQFOQQFQON```````````````````
(�B� @�	�&L�2dΝ:t�ӧN�:t�ӧR�J�*T�R�J�*T�R�J�Jdɓ&L�2dɗ.\�r�˗.\�r�˗.L�Je˖�Z�jիV�Z�jիGq�q�q�q֭Z�jիGq�q�q�qݻv�۷n�qݭL��S�I�J�)5#�L�2R�ҕ )4���R�JR�S��R�� �T�\�2��
��'I�L� ��$ʣ!�������@Kӎ�O1/C
�d��@S���D0AuAabW�s���/Qb��)D��D(S���D5� "&H���3n���,"���]	&ǆȧ��*�B�#O�щqy钊��q���2p�p��r2���)q(���(��s���{����n7 ����q��o�q��I� �~���A�o`������� ]d������%.%%%.../////////12FQQQQOOQQQON`
(P�B�
(P�B�
(�D @�*T�R�J�:t�ӧN�:t�ӧN�J�*T�R�J�*T�R�J�J�ɓ&\�r�˗.\�r�˗.bŋ,X�b�2�)�1Z�jիV�q�q�q�q�q�q�Z�jիV�q�q�q�q�v�۷nݻq�,:�)R�Lt�f*J��\�j�+�&Rt�S�S&\Ŋ��R�J�r�ɔ�Z�k�N�JT�2�T�R�*d�J���2�zqꠠ�!��&�J�(�(�3�T�*��M�D���r2����*T���N�:��0�O@d��Z{�E��}��<�d	����/�'3Sb""�I�XC�]y%��%��YX����u���***!�����QC=T.%221C1%=/=%.12/=%�������8�`� �78� 8����?��7��3��,����������������**��*(����������0
(P�B�(P�B�
(Qɓ&L�2dɕ*T�R�J�J�*T�R�J�*T�R�J�*T�R�J�*T�R�R�Jd˗.\�r�˗.\�r�˗1bŋ,X�\�2d˘�Z�jիV�8�8�v�۷nݎ8�8�Z�jիV�8�8�v�۷nݻv�۷nݎ8�v�2�)�)R�j�jF.bŊգ��2�*T�LŊիX�L���˘��۷c�L��aئR����N�R�)T�T�QF`FTQ&�2ypr3U)��Q`@��S*�A�T�B�:T��������
u)2�(�NTQ=u�Ӟ�f���&U*1s��H�|����2�$>^k�M��J���-���RRUC# ���K�(���*!�����#�������������������b�XK��� q��:��7�@�".�%./u���OK�E���K�OOK���LOK�P̑�TOLP��TTS�TQ�SӘ @�
@�2dɓ&L�2dʕ*T�R�R�J�*T�R�J�*T�T�R�J�*T�R�J�*T�R�2e˗.\�r�˘�bŋ,X�bŋ,X�\�2�,Gq�q�q�qݻv�۷n�q�q֭Z�jիGq�qݻv�۷nݻv�۷n�qݎ���+V��r�+���۷nݻv�u�W.b�q֭Zŋ�q�u�GwnݭZ�jիV�b�r�ɓ)R��2�'&t���d�IS%*L�T�R�J�*T�R�J�*T�N�:T�R�J�*T�T�N�*T� @�yHg�F!��ʰ
u��������v��҃8��i"��
!IrHJ�S#�deEDde����edeEEEC##$443������rRR�Qq`��Hc��    �u���:� η��)qq)(����))yyy����������������222���222��zzzrrs P��(Q	� @�2eJ�*T�R�J�*T�R�J�J�*T�R�R�*U+��J�*T�R�J�*T�R�L�2dɓ.\�r�˗.\�r�˗1bŋ,X�bŊիGq�q�q�q�v�۷nݻv�۱�Z�jիV�Z�q�q�۷nݻv�q�v�bŋ,Y��X�Z���)�1Z�۷nݻv���X�\�h�Z��#�8�8�V�8�v�jիV�Zŋ˓&L�J��I� �T�N�
�e�J�&�*T�R�J�*T�R�J�*S�N�*t�ӧN�:t�ӧN�:L�2dɓ&A)UD��2�
'E�/ ���3�˓JH���..�n��@�������U��Q��S�ӓ����TTTTTQ��������LLLK��OOIK��K�Eş�!!���!!!!  /���$1��  ��ˏOOK�E��K�K��LLP����������̌�������TQ�����ӓ���(P�B� L�ɓ*T�R�J�*T�ӧN�:t�T�R�J�*�)R�R��T�R�J�*T�R�J�*dɓ&L�2�˗.\�r�˗.\�s,X�bŊ�,X�Z�q�q�q�q�wnݻv�۷nݻu�V�Z�jիGq�qݻv�۷n�wn�,X�bŝ�u�V�k+Gv�۷nݻv�u�W.b�q�Z�k#�8�8�8�8�V�Z�jլX�\�rd˗&Rt�2aHL�r��T�b��2iR�J�*T�R�J�*T�R�Jt�ҧN�:t�ӧN�J�J�%J�*T�R�T�NOA�)43$�.� �Tg�����y�)
���Q+݀)�R
��ΰ'�`NOOOON`NNNNOOOQOQQQFFFFTTT22CCCC111////=//1/=.%{��BBB@@C�������Ã�����XK�X���ļ������������QQQEEE===EEE9999��(P�B�(QD&L�2dɓ*T�ҥJ�*T�S�N�:t�ԩR�J�*U*R�J�s*T�R�J�*T�R�J�˗.\�r�˗.\�r�˗.\�r�,X�bŋ�X�Z�h�8�8�8�8�ݻv�۷nݻv8�V�Z�jիV�8�8�v�۷nݎ8�ݖ,X�bŝ�v���V�v8��۷nݻv�۱ֱ\���c�:իX�8�8�8�V�Z�jիV�Z�j�,W.\��ɒ�*U�QU+��b���T�&UJ�*T�R�J�*T�R�J��R�:t�ӧN�:t�өT�L��ӧN�:t�QI�,�

bd�Pc�9��#�L%EP����X�OQ:)ԡX

����Srrrzzzzzz��2222��������yy���y�s���������IIK���Ń��w��X���ļ�����QQQQQQQQQEEE==999==EEE9���(P���(�&L�R�I�*T�өN�:t�ӧN�:t�ӧT�R�J�*T�J�*��T�R�J�*T�R�J�*W.\�r�˗.\�r�˗.\�r�˘�bŋ,W1b�jգ�8�8�8�8�v�۷nݻv���Z8�8�8�8��۷nݻv8�vX�bŋZ;���Z�۷e�;v�۷nݻv���X�\�k�n�jգ�8�8�:լX�Z�jիV�Z�k,W.Z�re)N�N`U*e�X�j��R�R�J�*T�R�J�*T�R�JT�N�J�*T�R�:u*T�T�J�*T�R� �99���y�11F%�AH'��	'����F&u�=8��d	�*�QB��(�P�X���������TTTQ��������LP̌���K�EŃ��p�aqqqrRR�����Qqa`縱)y�����������������222222222���zzzsrrrzz{ P�E
(Q	�&L�2�N�:T�ӧR�Jt�ӧN�:�*T�R�J�J�*T�R�JT�T�b�2dɓ&L�2dɓ&L�r�˗.\�r�˗.\�r�˗.\ŋ,X�b��+V�q�q�q�q�۷nݻv�۷n�j��q�q�q�wnݻv�۱�۲ŋ,X���;Z�J�ݖ,�u�ݻv�۷n�Z�r�+]�v�q֭q�q�v8�X�\�jիV�Z�u�V�b�s+�):t� RT�\�j�*N�L�J�*T�R�J�*T�R�2�*R�J�*T�R�J�)ӧJ�*t�ӧN�:���ӓ£(���00O*<� �����b��0
 @PRB�:T�P���(��

+rrzzz����222��������������q(��������)))qqqy��q(�����q�������������222����������zzrrrpV����B�@�&T�R�J�:u*S�N�J�J��N�:t�ԩR�J�*U*T�R�J�*R�J�sɓ&L�2dɓ&L�2f,X�bŋ˗.\�r�˗.\�r�,X�bŋ�X�Z�h�8�8�8�8�ݻv�۷nݻv8�V�8�8�8�8�v�۷nݎ8�ݖ,X�bœ.۵���Z�gkX�v�۷nݻk˘�,Y۱�q�q�wn�Z�re+V�Z�jգ��j�,X�\�JS�I�@�T��&\�2T���L�2dɓ&L�2dɓ&L�J��R�J�*T�R�R��1AB�:t�ӧN�`
��1y���B�R�Q&AQ��2��N:t�2d
�:�UI�	�&@PP��(P��X�00''''������###***!�***����������������������������*!����****###(�������������''00
���98P�B�&L�2dʕ*t�S�R�J�*T�T�L�*T�R�J�*T�R�J�2dɓ&L�J��R�\�2dɓ&L�2dɓ&L��,X�b�r�˗.\�r�˗.\��,X�b�s,V�Z8�8�8�8�;�nݻv�۷nݎ:ծݻv�۷c�8�8�ݻv�۷c�;�e�,X�d��������,Y���ݻv�۷n�Z�r�+Kv���8�8����W&R�jիV�Z�q֭Zŋ˓):T�2�I�:�s�S)J�p�&L�2dɓ&L�2dɓ&R�JT�T�R�J�)�%*A�9<�R�J�*U9QD��׸��H���E(�&:�)�92��!R�
R���T�SήJ@�T�

Q
((P�B�00''''������###***!�**!�����������������������������!�!����***###(�������������''000

+p�B�&L�2dʕ*t�ӧR�J�JT�T�L�2T�R�J�*�*T�R�Jdɓ&L�2�)R�R��dɓ&L�2dɓ&L�3,X�bŊ�˗.\�r�˗.\�s,X�bŊ�,X�Z�q�q�q�q�wnݻv�۷nݻu�]�v�۷n�q�qݻv�۷n�wn�,X�bîR���\ň���۱�j�n�jիV�Z8�ݻ,X�bŋjլX�b�3ݻv�۱�jլW&Jt�Dɕ*T�ӣ�Z�rd�T�R�J�*R�R�JS�R�J��ӥR�R�2�,R�*LSrqB�
���dd��P�P��X��� (Qdʕ:t�T�R�J�*T�T�R�*S�I�&@�B�� ((VB�
(P����dc###%EEDc#######"�����������443��������4444dddddddeEEDde��������X����
(P�B�
(P�B��*T�ӧR�R�Jdɓ&L�2dɒ�J��ӥS&L�2dɓ&L�2dɗ):u3ɓ&L�2dɗ.\�r�˗.\�r�˖�b�r�˓&L�2dɔ�L�2�ˇq�qرbŋ,X�bŋ,W.\�r�˗1b�jի]�v�۷n�,X�bŋ,Y۷c�0`��0`딦b8�X�Z;��%�;v�q�v��㎵j��۷n�q�q�u�V�b�3ݻv�۱�jլX�R��2	�&L�s+�&R�)ӫ�.\�r�ɗ1b�2���.L�2�$ɕ*u*U)N�&(*rrT�R�J�+���Rd�0@�S��
(Qdʕ*t�ԧN�:t�өR�:t�R�J�&L�

������������������������������������dd���bbb^^^^bbbbzzzz^^^b����dd��������������������������(PP�X�
(P�H @�&L�R�N�:�*U*R�J�*T�T�J�)ӧS&L�2dɓ&L�2dɗ):u2�ɓ&L�2dɗ.\�r�˗.\�r�˖�b�r�ɗ.\�r�˓&L�r�,V�Z�jիX�bŋ,X�bŋ,X�bŋ,X�b�j��v�۷nݻ,X�bŋ,X��n�`��0`��b�2��Z�qݖ2X�b�ݻ�gnݎ8�;�n�q�q�v��㎵je�Gv���ݎ8�V�Z���)N�bŋ�V��qֱb�r�˗.\�re˗.L�+˗&L�J�*S&\�r�ɒ�*L� P�E
)Dļ�E�)2d�(Q2d
 L�R�J�:�)R�J�*T�ӧJ�*L�R�J�&L��AB�''��00000000'''��#***###(�����������*!��������������������***###(����������������
(P�B� @��B��
(P�B�&L�2dɐ&L�R�J�*T�өR�:t�ӧN�R�JT�R�L�2dɓ)R�J�*T�Rt�˓.\�r�˗.\�r�˗.\�r�˗1b�r�ɓ1bŋ,X�\��+V�Z�jիV�bŋ,X�bŋ,X�Z�jիV�Z�h��q�q��bŋ,X�b�ݎ8�,X�bŋ,;˖�v8�vX`��,Y۷e�v���8�vX��nݻv��b�ݻq�.Z;��Z��㎵j�֭b�2�)�&L�s.ݎ��˔�R�J�*R�R�JR�S)R�*T�T�R�2dɔ�Jt�2�:�Jdɘ����P�B� @�ӥI�*t�өR�R�IӧN�:t�T�N�:T�ӥJ�&L�2```
(P�B�
��9=EE���QQQQ�����QP��������QQEEE==========EE===998P�B�
(�2d�(� @�R�J�*T�R�N�J��ӧR�J�*T�R�J�2e*T�J�2dɓ&L�J�*T�R�rR�T�\�r�˗.\�r�˗.\�r�˗.\��˗&L��,X�b�s,V�Z�jիV�Z��,X�bŋ,X�b�q�q�jգ�;�c�8�8�ݻv�۷e��v8��۷nݻv�۷n֮\�۱ݻv��bŋ,Y۱�,Y۱�u�V�8�ݖ,X�bŋ,�۱�s��:ծݎ8�V�u�X�\�2dɗ.b�rd�R�:Ur�˗.\�*�ɔ�:U2e*T�J��2d @�2d

�2�N�:t(P���)����HL�j�)N�J�J�*S&\�r�*T�R�Jd�T�J�)R�J�&@�ҥI�(P�B�
(Q��0''**##(������������##***'���#*****###(���##(������������������''
(P�B�&L�B�&L�2dɓ&L�2dɝ:u*T�T�J�*�*S)R�J�*T�R�JT�N�R�J�*T�R�J�*T�JT��ɔ�\�r�˗.\�r�˗.\�r�˗.\�rdɔ�bŋ,X�bŊիV�bŋ,X�bŋ,X�bŋ,X�8�8�Z�h�8�8�;�nݻv�۷n�u�]�v�۷nݻv���ˇ,�q�q�wnݎ8�V�v8�V�Z��+V�ZX�bŋ,�۱�j�+Gqֱv�q�Z�jիX�b�s,X�Z�wc����ɘ�bŋ,S&\�re)S&L�J��T�J��ӥW.L�2�*I�&@�B�*L���J�&L�
R�:t�U)R�R�2d�R�J�*T���R�*S�ɓ @��GJ�&@��B�
(P�B�`NNOONNN```
��������999===EE=EEP��QQQEEEQQQQE========EEEE===999999998P�AB�``(P�B�
(P�B�
&T�S�N�:t�T�T�R�J�*T�J�*S�J�J�*T�R�J�*T�R�Lt�T��)L�2dɓ&\�r�˗.\�r�˗.\�rd�T�bŋ,X�\�s,V�bŋ,X�bŋ,X�bŋ,X�Z�jիV�\���V�Z�jիV�q�q�v�q�Z�h�8�8�9e���X���Z�j�,Gu�X�b�jլX�\�2e˗1b�jիV�Z8�Z���Gu�W;v8�Z��,X�b�2dɗ.b���b�re*T�R�J��N�:T�d� (P�*R�:T�3�N�*T�T�R�&@PR�I�**0FFFTTT22*L��D	� L�2�J�*T�R�J�:t�R�ɓ @��AB� @���	�����������*(ʊ�H��*)��������������ʊ��FJ��Hf%��&&(hfFFHhhhfFJ��*******(����*)����������	���������������������B�
(Q&L�R�J�*T�R�N�*T�2eJ�*T�R�R�J�*T�N�*�2e*T�R�J�+�.\�r�˗.\�r�˗&L�J�+�.\�r�ɓ&\�s,X�bŋ,X�bŋ,X�bŋ,X�bŋ)�.\��+V�Z�jգ�8�8��u�V�Z�jիV�Z�j��W1�gkV�bŊ��V�bŊ��X�b�r��T�L�2�˗.\�r�íZ��,V�8�b�۱�jի�1bŋ$ɕ*T�Ӣ��`NNOO
(P�B�OONNNOQFFFFTTT22FFT2CC11	u��_�0g������H�%T` +rs P�B�(P�B�
(Q
(�B��
��+rzz��������������yyyyyy��qqqqqqqq���qq)))��y�(���qqq��yyyyy��22222222���22�����������rzzz������������zzzzzzzz��zzzrrs P�E
(P�B�
T�R�ɐ T�R�J�*�*T�R�J��2iS)J�*T�R�J�r�˗.\�r�˗.\�2d�T�R�2dɓ&L�Jdɗ.\�r�˗.\ŋ,X�bŋ,X�b�r�˗.\�Jd˗.\�jիV�Z8�8�8㎵k+V�Z�jիV�Z�ƙE52�*T�R�JT�R�J�*��R�*L�Rd�

�E9�=P���������\8$�^.�$u�� :� IP̋����������ѐ�E�]` /p����%�.z^zJ,�u���:�b0pw����~�^o0ppw���q��n0w�#�h!��t<��"�(����������������	������***(��ʈf&(j��%ʈg���������������秧����ǥ����(j��w�qyqrz�����y���b����[��������?��2��*#(�00(��'�

�����dbz\���������Q�2r2��������zzzzzzzzrrrrrrrp�B�
(Q2dɓ&L�R�J�*T�ӧR�J�JT�T�L�2�˗.\�rdɓ&L�2dɓ&L�2�˗.\�r�)N�J�Jdɓ&L�2dɓ&L�2�˗.\�s,X�bŊbhǢ��$	�R�k��ݻv�۷nݻv�۷e�,X�bŋ- Lv)R�*T�R�J�:t�ӧN�NNOQFT2C%%%%?�������/T/%	WX3u ��=ˌ��EŅ��US��B�'�����###*���#������������**!�00
(�ddddddde�$543%Dde�B�
(QB� L�0�B�0'''
((V��єTQ�NF22TFFFFFFFFFTT22CCCC./=%%..%%=/%%u���@	�7H����u�_�1arR���5��P�
(Q0'�
 8(�(�D	�*U<�Rd	�&L�2dɓ&L�2dɓ:t�ӧN�*T�R�J�*T�R�J�*T�R�J�:t�T�T�J�J�ɓ&\�r�˗.L�2dɓ&L�2dɓ&L�2dɓ&Z����V�\�r�˗.\�r�˗.\�r�˗.bŋ,X�Z��V �ΩR����v�۷nݻv�۷nݻ,X�bŋ,X�a�&*t�R�J�*T�2dɓ&L�P�	��*"�
������(�B�`NON
@����ST�QK�H'�RŊc�N�
��Rb�� 9EPP�eJ�&M=8(�L
(�E

��T�2d
��������L�2dɓ&���=EE<�Rd`N(P�B�
&L�R�N� @��B��&L�
*�QE98�T�dddddddddddc#$443R�42����W�ܸ��X\�X�8���2	u��I���AFJ�K��OK�P���X�
dJ��������@P�AB�`QO`@�2lB�(P�ΥR�J�*T�R�J�*T�R�r�˗.\�J�*T�R��ӧN�:u*T�R�J��ԩR�R�*U*S&L�r�˗.\�r�˗.\�r�˗.\�2dɓ&L�k˗.b�r�˗.\�r�˗.\��,X�b�jիV�Z�j�,V�-wn�,1۷nݻv�۷nݻv�bŋ,X�bł�v�8��R�J�*T�I�&L�2dԥJt�R�H @�B��`2/2`:��2ԭ,��T��.�-LŊ�gR�JT���:��S�N�&L�ʝJt�R�N�*@+ �D	� (S�
(SS������ L�T��������D&L�R�J�&L�
(QI�)�I� +z���2��������zz���222221��2p�l
���*'��������ӔH1QQ%QO=.QOONN``
�1(�z�rzrs P��F ��r��,�:t��dɓ&L�6&N��D�S��:t�ӧN�:t�ӧT�R�J�*T�R�J�*T�R�J�*T�R�J�*N�J�J�)��R�2dɗ.\�r�˗.\�r�˗.\�r�˔�R�J�*R�*T�S�X�bŋ,X�bŋ,V�Z�jիV�Z�jիS.Z�bņ,Y۷nݻv�۷nݻv�۷n�,X�bŋ,Ys�H%ZL�R�J�*T�R�J�*T�Rdɓ&LP�B�
)jT�wX Hsz2�34�ҦL�I�ʅ`&t�ӥN�:L��d	�Jt�ӧN�J�)eN�:T��)R�*@��ʕ&@Q2dɓ&T�T�N�*T� @�b�ʈ�)ʈ�)�H:��������L�2�J�:�*S�J�*T�2d� t�T˔�O*T�Rd
&L�2dɓ*T�2dNO2=%/Q���{�?��LD���j�!��!!�1 �� ����}>�BBBBD�G\�^���QE8(�0�C����2��2����������W���P�b�J�*T�R�J�*T�T�R�J�*T�R�J�*Tɓ&L�2dɓ&L�2d�R�R�2d�T�L�2e˗.\�r�˗.\�r�˗.\�r�ɓ&L�2b�I� L�U�V�Z�jիV�Z�j��q�q�q�u�Gv�v+�v8�V�v�۷nݻv�۷nݻ,X�bŋ,X�e!��lJ�R@� �*T�R�Jt�ӧN�:�r�,V�Z��$�JS�S-QU��;b�h�e����Z�rլS&@�ԧI�J�*T�R�:�Jd�R�R��ӧN�:�J��N�:u*U*T�&@PP�J�*T�R�LOP��``
P�D	�&L�2dҩR�2d˔�J�)ӧS&R�JT�N�J��y(HQD��@� ����������b.Jd���*\z�^?�,�G�N"!B��gp}�@�*|Y��"�|��&b�Y�1f,Ř�dm����.^b�d�����)8�YP� P�X��(PP�B�
������*T�R�J�*T�R�J�2dɓ&Lt�ӧN�:�2dɓ&L�2dɓ&L�*�)�&L�*�)�&L�r�˗.\ŋ,X�bŋ,X�b�r�˗.\�2��T�\8�8�8�8�8�8��۷nݻv��b��b�q�Z��.ݻv�۷nݻv�۷e�,X�bŋ,@+�S:t�ӧN�L�2dɓ.\�s,X�*T�T�T�:�j��L�2dɓ&v��T��	��\�ie�T�
�RN�&U*��S&L�J�*R�L�r�ɔ�J�*�˔�L�rd�I�*t�T�GZ�re)R� @�)&��U2�
(P�EJ�*T�R�T�R�2d�T�J��ө�&R�*T��
�d.���+z2rrrrrrrr�������22��� �į5fAf�p'�>NGDR}ȊO��N �'f�G��f%4�3L�2̳,��>'	���2z���22���)N�*L� QDʕ*L�Rd�
))ԥH*�*T�R�J�*T�R�J�2dɓ&L�*T�R�J�J�*T�R�2dɓ&L�J�)�.\�*�)�&L�r�˗.\ŋ,X�bŋ,X�bŋ,X�b8�X�Z8�8�8�8�8�ݻv�۷nݻv�۷e�;v�q�q�q�v�۷nݻv�۷nݻ,X�bŋ,X�j�e��bTq�q��,X�b�*U*T�L�J�˘�Z�v�����1Z:�ɔ�R�re+rɉ�Z�ltɇ,:�'J�R�JV,W.L�J��T�\�2�)R�R�h�T�\�2��R�R�r�)��:T�GN�:t�Ӥ§�
�b����Qb�
(P�Dɓ*T�ӪT�J��ӧN�*T�2gI�*�I�d	�R��2 @�
((P�I�Γ
���ļ���!0GX` ;���{�?_�1�@@��0XRrrrzzz���b�X c��$�{:�N�P0i�����}�����g�k�I�buh�ɓ&L�2eJ�*T�R�N�:t�ө�&L�2d�T�R�J�)�&L�2d�T�L�2��R�R�2d˗.\�r��X�bŋ,X�bŋ+V�Z�jգ������۷nݻv�۷nݻv�۷nݻvX�bŋ,:�,X�����b��v�۷nݻv�۷n�,X�bŋ,Y��Gv:�]���;v�۷nݻv�۷nݭZŋ��q�q�v�۷nݻZ����V�q�q����V�R@�S�I�R�s�c�\�2dɗ.b�r�˗.\�r�˗.\�J�)�.\�*T�R�J��R�R�R��dԝ
���r�y4�I�T���ɔB�����eHLtɒ�*M=*��J�&u)�
&E礤�����������������·����~�>�@�"���� G����J�q������ N���%g&��VV�F�A�8,��P�a�zj�2c��D"ٖi�~C��A��D��O����2�t	�&�*T�R�J�J�*T�R�L�2dɓ&R�J�*T�R�J�*T�L�2dɓ&\�r�˗.L�2dɓ&L�r��X�bŋ,X�bŋ,X�Z�jիV�Z�jիV�Z�h����8�;�nݻv��bŋ,X��8�;�nݻv�۷nݻv��bŋ,X�bŋ,X�bŋ;Z�h�W%Z���X�Y۷nݻv�۷nݻv�j�,X���8�;�nݻv��լW.b�h�8�8�W.Z�r�R�*Lꓩ���2�ɓ&L�s+�.\�r�˗.\�r��T�L�r��T�R�J�%N�J�Jd˗%J�1Ri�T�NuH��	��# )J��q4�R����3�S.J��T7���H�ڲ�ʪ����������ffffffff�y<��.��g���H�}��o�؈��D5��#���$@�|>ܳM�Ӆ��p��:���` ������.�=2.��������������   8�N��R�J�*T�T�R�J�*dɓ&L�2�*T�R�J�*T�R�Jdɓ&L�2�˗.\�rdɓ&L�2d˗.bŋ,X�bŋ,X�bŊիV�Z�jիV�Z�jիGwn�q�qݻv�۷n�,X�bŇq�qݻv�۷nݻv�۷n�,X�bŋ,X�bŋ,Xv)�1Z�*�n�b�r�ݻv�۷nݻv�۷kV�b�h��q�qݻv�۷n�Z�r�+Gq�q����V�RLꔥI�Ru3)��L�2d˗1b�r�˗.\�r�˗.\�J�ɗ.\�2dɓ&L�*�*S&L�2�˓% M2baH*�\J���p���^�H�)*a��H
*�re)�I�&L꒥N�J�2gnݻv�ۿ�����6�l��q���hL�Mo
>3�ņ;v�۱�����%J�r��N�:t�өR�J�*T�T�R�J�*T�R�J�*T�R�J�)�&L�2d˗.\�r�ɓ&L�2dɓ.\��,X�bŋ,X�bŋ+V�Z�jիV�Z�jիV�qݻq�q�v�۷nݻ,X�bŋq�q�v�۷nݻv�۷nݻ,X�bŋ,X�bŋ,X�e���\�r��ݎň坻v�۷nݻv�۷n֭bŊ�ݎ8�8�v�۷nݎ��,V�8�8�;˖�\��U)J�*�J�W)L�2dɗ.b�r�˗.\�r�˗.\�J�)�.\�r�˗.\�Jdɓ&L�qT���J*����&��2 ��|�՜ ��`*���Ri�N�L�+q+]���a��۷nݻv�۷nݻv�Jd�V��۱�u�V���Y1#����̆����1gc�,:�+��,Y�a��n�\�q�ݎ����X�b�r�ˣ}*T�R�J�*T�R�J�J�*T�R�J�*T�R�J�*T�R�2dɓ&L�r�˗.\�2dɓ&L�2e˗1bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�jգ�;�c�8�8�ݻv�۷e�,X�bÎ8�8�ݻv�۷nݻv�۷e�,X�bŋ,X�bŋ,�rT���\�۱ر��nݻv�۷nݻv��լX�Z;��q�wnݻv�۱�ZŊ��q�q����V�R�Je%I�J�h�W.b:dɓ.\Ŋ�˗.\�r�˗.\�r�*S&\�r�˗.\�rdɓ&L�J�jV�R��JRԥ
^H�/T{����$���:ь�T�	���d�:�S�]��h�ݻv�۷nݻv�۷nݻv�۷���;Z�30|�8%�XMZА��F�u*j]�0gb�JS�R�Z�*T�W&\�r�˗.L�r�˗. MK!S�%J�*T�R�J�*T�R�R�J�*T�R�J�*T�R�J�*T�L�2dɓ.\�r�˗&L�2dɓ&L�r�,X�bŋ,X�bŋ,X�Z�jիV�Z�jիV�Z�q�v�q�q�۷nݻv�bŋ,Xq�q�۷nݻv�۷nݻv�bŋ,X�bŋ,X�bŇ\�*e���۱ر��nݻv�۷nݻv��լX�Z;��q�wnݻv�۷c�Z�h��q�q�b�rի��L�1�eN�Z��d�]�L�2��X�\�r�˗.\�r�˗)R�2e˗.\�r�˗&L�J�)R� ��U#� ��u���b��0�+���)H;�}�$&�7X3)C�=:��yņrŝ�k,X�bŋ+V�Z�jթ�)R�*T��\�� ��	�&E���ϣr���Å����!����zdL��ļ]��=NOFT2222�^��=99�(�D
P�
@�1G]�:t�ӧN�J�*T�R�J�*T�R�R�J�*T�R�J�*T�L�2dɓ.\�r�˗&L�2dɓ&L�r�,X�bŋ,X�bŋ,X�Z�jիV�Z�jիV�Z�q�v�q�q�۷nݻv�bŋ,Xq�q�۷nݻv�۷nݻv�bŋ,X�bŋ,X�bŝ�J�0�-v�v,G,�۷nݻv�۷nݻv�k,V��q�q�۷nݻv���Z8��q�q�b�rի��\�1�eN�\�)ө��L�2��X�\�r�˗.\�r�˗)R�2e˗&L�2dɓ&L�JS�J�Q*�<�c$cS�C�
�p��D��M�-I+
�"F�U�vՃ��A�`���,�<�R
*$ (P�I����������������	����(����e��w����y�2���b�0������ �  ����*���0'��#(��0
OTTN
���(QB�
(Qdʕ袩N�LT�R�J�*�*T�R�J�*T�R�J�J�*T�R�J�*T�R�2dɓ&L�r�˗.\�2dɓ&L�2�˘�bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�j��۱�q�wnݻv�۲ŋ,X�a�q�wnݻv�۷nݻv�۲ŋ,X�bŋ,X�bŋ,�JUÌ�۱ر��nݻv�۷nݻv��լX�Z;��q�wnݻv�۷n�Z�wn�q�q�b�rի��b�1�dΥJ���	W&L�2��X�\�r�˗.\�r�˗)R�2e˗&L�2dɓ&R�)ҥI�%Q z�(X8%����0#t4̒���Ԫ��f�6<7GD4Xa?<�h��/�r�@�N� @���QQE========P��ļ�]��{�����=��3F�f��ϋ{{	��lh�6�ގ�O	2.%{�Ë��OOK�ѓ�
��Q �B�'''��
(�2eL_�&IW
T�R�J�*�*T�R�J�*T�R�J�J�*T�R�J�*T�R�2dɓ&L�r�˗.\�2dɓ&L�2�˘�bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�j��۱�q�wnݻv�۲ŋ,X�a�q�wnݻv�۷nݻv�۲ŋ,X�bŋ,X�bŋ,��˖�0��X�X`�kX�Z�`�8�;�֭Z�we��k+��Z�jիF;Z9a��b�wn�Z��d�G\�2��I�(��H(��bU2�ҦLT�T˗&L�IQD�&*�*r�!a�&b�)+N�J�t�礠!��o���0@wؑ�fS�i���Ъؾ��h��<4GGGggggBp�M�Z/78�z�����g�I��J���.@��2z�qOr�����BOS˟η��8�%QƢ�12r?� ����l6�h�hx�Ԫ����JLXX�=����OSÉJ�!�����'& �����^�@�VgI�{��
:t�JS�I�*t�ӧN�:u*T�R�J��ԪT�\�J�*T�R�2dɓ&L�J�*T�R�2dɓ&L�2dɗ.bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�q�q�q�q�q�q�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�bŋ,X�bŋ;Z�s��v;+]�,:�˖�Y۱�q�u�X�wn�k+�q�q��r��b�q�k˔�reɔ�*@+pRª*
RU2�b��:T�Tɓ&R��q���b��!�% �2���S�S��J� ,\  �}8\.��g	���SkC*�B�J��H���""Z�P�"K����u��	��� M<����3aI�TJ�
`=F2OQ/%/CC%/OQ���\o���s�y�8���3��0kAD<WXGYFO���
2Cu���?�OKß�JTS���O
��@PQDΥ
T�U��N�&L�R�J�*T�R�R�J�*T�N�J�2d�T�R�J�)�&L�2d�T�R�J�)�&L�2dɓ&L�s,X�bŋ,X�bŋ+V�Z�jիV�Z�jգ�8�8�8�8�8�8�ݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷e�,X�bŋ,�u�X��gc�b�q�Z�r�+Gv�۱�u�W.\���n�ZŊ��V�Z�jծ�b��aֱbŋ,X�L����S%J��6c%44�eS) ���D (�T0�d5C�c��P�SӉE����=u���_�7P;�i��s	��ښ�ZZ[[[[U�YOL�NNNNU����[�І���" ��w	s�Ɯ�D�0�a'� ��**�� %���ǥ����eΰ��c�����' �$y�3,�B�2׍�F���M��.r�w��� \��.	{��������'�!�Q1�QRl��J���6%J� @�eJ�*T�R�N�:t�ӧN�:�*�*T�R�J�*T�R�J�*T�R�J�*S&L�2dɓ&L�r�,X�bŋ,X�bŋ,V�Z�jիV�Z�jիGq�q�q�q�q�qݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷n�,X�bŋ,YjիV�;�n�Zŋ+�.L�r��ݎ:լX�L�J�)��kɓ)L�2dɓ&���GZ�rd�T�L�qR	T�&T�S�H'���##��'�Ju�E9D������9D���%=�� �:�������_䪈opG���}����7L۠o'�'''''����Ɔ���օUT��������C�q�cE���ɛ[�5a�&�t���\�.bR���bQu@�&%��ʆ! &D�&G�w�s�]�ͷ/�GG�|��!�,>~#
,� ���QC�'��:Kk��}��&H`)�j��'�qvc1e�)��'��0(�J@PP�E&@� T�R�J�*t�ӧR�J�*T�R�J�J�*T�R�J�*T�R�2dɓ&L�2d˗1bŋ,X�bŋ,X�b�jիV�Z�jիV�Z8�8�8�8�8�8��۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻvX�bŋ,X�b˗1Z�q�qֱ\�J�*S&R�H�X�\�J�)N�:u*�+�&R�)�dɓ&L�5ɒ�\�2U)N�*u*��	�0'0L�US442��3&d�̕�K��OK�E�P�E�˅� C�qg�	��Q�8��{���=�`���#���y8].wK���|���L������\��W�YYYUURRRW�W�W�QNU�� �O�apg;cHC{c�� bd �=u��*F==O%u���?IS�\��=f�>��"�afbE����H58���$T���#!$��� ��}y��y=�g���fE�*�fL	ʈ��)���(i�TP�`O:�����QB�
(P� @��N�*T�T�R�J�*U*T�R�J�*T�R�J�ɓ&L�2dɓ&\��,X�bŋ,X�bŋ�V�Z�jիV�Z�j��q�q�q�q�q�wnݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۲ŋ,X�bŋ:�3�X�Z8�X�Jt�ԪT�:Ure)N�&@�Rdɓ*uJ��J�&L(P�B�
)�eR�:L�1L��
�d�����������bzbbbbbbbb����zb�bz^^b^z\J.zzJ\z �	����ˌ^�Xp`�� �}�@���@�-���Cu��3VzjirxzVxhYxhhhh__eeYIXleIle_4@W@D9<<z@^ir<WGgWk<lHn�2���/���R��X���.�t ����I&��.4ܑ����?�� ��!"6�8����%4��B,��d[r֐�D_}>�"b�IA� "��S§��*M1T�kJ��OOQOO`@(P�B�
P�B�
(�ҥI�&A*T�R�J�*T�R�J�J�*T�R�2dɓ&L�2dɗ.bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�q�q�q�q�q�q�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�bŋ,X�bŉ�R��ɖ�v*N� T�'J�Jt�1AS��� (QdΕ*L��AX
�(�Rb�OQQO
A�QE=P�QEQP�����������QP���ļ��ļ��\X�]�,\.\�.	�����w�pH#�A��{	�@�N00!��K�!��s��++�+((=<5554������4/����*����+�$��#���3��"$�"��#��� �2��5��:JUYP���C���\H��Q�m��qۀ� ��q$#��/�$�	>'����Q8\h���&|Y�Q�B��A���o��b�@FAR�NFFFFQN
)��������(P�B�
�Ҥɐ (�ӧN�:u*T�R�J�J�*T�R�2dɓ&L�2dɗ.bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�q�q�q�q�q�q�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�bŋ,X�bŅJ���X�v*J�L�T�I�*L�V�bd
(�2d�
��(P�B�
�V �
`��dd��(*���r1�22��2������*p���)qqq(�s�\]��	%1=u��������@@��u���bn�0�'H��	��t�F���.NwɛÓ�������K�Cj�ª��B#cj���+*JJ�+cA���:I��b;CC9�"
ª�"��t��x̑�bPőW��QZY�|�j�D(���ř#0��� ��͙VJ/��E���ςq~[��B}��g��,.'I�P�)&��⼲f�f�mQ=ΝFTTTFQN
)��������(P�B�
�Ҥ�(�ӧN�:u*T�R�J�J�*T�R�2dɓ&L�2dɗ.bŋ,X�bŋ,X�b�jիV�Z�jիV�Z�q�q�q�q�q�q�۷nݻv�۷nݻv�۷nݻv�۷nݻv�۷nݻv�bŋ,X�bŘ:��1GT�Z�1R��
������������(�B� @��B��
��QB��00''''��������������**'���!��������������������� � �~����qaqp��K���$}���o�����}��O�7�k�5��t�>_-�3���33PPVrzzrrrzxjjiYYYhhh__UUUeee__U_hheIIUUlI_elIYYelUirziE8*Ɉ��|}f.}��Y�������f�1�>!�pQHAXU@9lA?������|��#?-�|ͳ �Sr����h�l�Dp_AŹa8��#���/�G��R�n���?�J�'?ب�* �T���ŀ����i�'(ӈ&T�U)��R�J�*S&L�2dɓ&L�r�,S&\�s,X�bŋ,Gq�q�q�q�q�q�q�q�q�q�q�q�q�qݻv�۷nݻv�۷n֭wnݻv�۷nݻq�`
L�Ҥ:�r�'I�(PP�X�
(P�B�(Q
((V� ��
����99==EEEEEEEE99=EQQEQQP�EP�ļ��ļ�����XX\\����������\8X�XX]�z,,�	u��n�@3�I�""�}>�O����$�}��������\ O'K�hh!��n���g3��Rf��������������������в���������ʒ�f��Ҡ��r���t�?%�Y#6�'���A!B��!��>G�~#��-�f���?���6*��� +��盤��8�����q">!��ܾ$`�paq��������AN&���Ԇd�Fr$kYgBxVB~�Χ./
�\�������R�*z�)z��S.\�JT�N�R�J�*T�L�2dɓ&L�2��X�L�r�,X�bŋ,X�Z�jիV�Z�jիV�8�8�8�8�8�8�8�8�8�8�v�۷nݻv�۷nݭZ8�ݻv�۷nݻv8��Q2d

@��*N�&L�B�

(P�B�
P�D((P�	��E
(P�	������������	���(�ʉ���(ʆHfFHf%�秦%��秧��䤤���ǥ���he�Ǩoq 7�x�pH ;���HH�u		>�BBBBBBBBN�P���""&�{���@��O'K�h !�4�n���b�35g''�g'''����������������'������ �������6���pN������H��f�����h������H7E4DWII9WUmYXAmoO:�8.|8�Y���"ߐS�8�C�3 �F?Y3!�?��[�Z���|Qn[��*����zz�}5:�E0Lb0�z�2c� �Uk��&R�)ҥT�R�J�*S&L�2dɓ&L�r�,S&\�s,X�bŋ,V�Z�jիV�Z�jիGq�q�q�q�q�q�q�q�q�qݻv�۷n�q�q֭wnݻv�۷nݻq�`
P�B�'0*u)ӥJ�&@�B�
(P�B�(�B�``NNNON`
(PV �B�0''''��������0''���#''(���������������������������*!���(�8DE�_��'����u:�D��S���u:�D���P����""&&�{�����@�O'K���|�[�g3��Rf��������������䬬�����f�s��L�OJT
�8�|_�J�|���TW/,�r�D5a55?���C�y�)�"�cj������:#�D��f�Y��������>P�H�B� �F�Y�AĢq?������'���y>�78����YŹn�O&��V���\���)�!��3�#�`` �)ɕ*t�T�R�J�*dɓ&L�2dɓ.\Ŋd˗.bŋ,X�bŊիV�Z�jիV�Z�jիV�Z�h�8�8�8�8�8�8�8�;�nݻv���8�:գ��۷nݻv�۷c�8�B�
Q	�H*t�R�I�&@��B�
(PP��
 @�rrrzzzs P�X
���999999999�99=EQEQ���\�����������ļ���������ĽQQ�P��XM�. �}��BO���I�HHHHHHHHHHHHHHHH�u:�O�����{����<�N�����@C��s9��fffj

��NJ��


'ɚ�Ku��t�>,Œ3g�n�/�|Cӄ����@���$�$7���#�,��$����(9��w3��ɨͥ)b���>�#���q�����8�XO�
��	��``q5?�F�\G���F"2�Dt#�4ͼ or~���=�Yە�%���*t�R�I�&�*T�R�J�J�*T�R�2d˗1b�2�˘�bŋ,X�bŋ,X�bŋ,X�b�jիV�Z8�8�8�8�8�8�8�8�8�8�8�8㎵h�v�۷nݻv���9AB�L�P��&T�R�ɓ @��B�
(PP��
 @�rrrrzzz��{ P�X

+rrrrrrrrzzz�2�����y�q(����������������������蹋�]��q�ĉ	��BN�S��$$�u									>�O�17���t�F�O'H�@C���s��JJL������JJ\�b���5���ܑg��Y��Y#1dτ=>.E'��qx
j�S��l�xn�����ʮh�h�ʲԬR���ʪ��ʎ�G��9�	#���dCg�	����j�jސ�`j��j6h�j�oa8����\G����0q8��`�@}��n��D�f���� �g3|N��h,	�W&R��2��J�*T�T�R�J�*S&L�r�,S&\�s,X�bŋ,X�bŋ,X�bŋ,V�Z�jիGq�q�q�q�q�q�q�q�q�q֭Z�jիV�wnݻv�۷nݻq�&@PP�
�&L��D	�&L�
(P�B�

P�DNNOOOQQQQON`
���(P��B�0''''''''(��#*!�������������****!���*****����?�n�a'S�����$�u:�N�!!!'S���u:�N�S������$$$$$$u		>�o�17�hk���p�<�.���������n�\�f�u��|�\�.gHue�#��|�!BE�g��,>�(�'��As	�LҠ���t�&��f��̷C���x�`�	y��l��rb1�^Kzd?	�C�2b� �!��m������������lݭ�!��ս���Fd8�[��X\O�!�5���� )�4$Ciq�"�&n������X*�zpQDʝ:t�ӧN�J�*T�R�L�2e˘�L�r��X�bŋ,X�bŋ,X�bŋ,X�bŋ,X�q�q�q�q�q�q�q�q�Z�jիV�Z�jիV�Z�qݻv�۷nݻv�q��1AE:��Rd
 L�2
(� @(QB� A9===EEEE=9�+p�B��
��������������d��bbb������ddd�����������ddddd������dbzz.�t?]���M��t?]��BGS�HI��u:�D����Ą���·C����$$�}>�b"bog�hk�	��t�^O'K�hhhh hhi��t�@�C\.e���_	�3G��Ϳ'�&>ȇ��<Өdb8����B-�8[��3$c��f\�D�`�6μ8��G���B�ק��p"*���t&�cv�e���ca�����cd�V�f�S��A��qdXPC�n	�qd8$C��`�R�U�S4�i"ƅ�@���ɦZt�ӧN�:�*T�R�J�2d˗1b�2�˘�bŋ,X�b�r�˗.\�r�˗.\ŋ,X�b8�8�8�8�8�8�8�8㎵jիV�Z�jիV�Z�h�v�۷nݻv���9ӥJ�&L�R�J�*T�2dɓ&L�2dɐ (Rs QB��''��������
(P�B�(PP�X���������TQ����TTTQ����S����TS�ё��TTU�̑��^�����u?D ���Ą��Ρ'P00����$�}>�_N�g���I�$�}�_�/�'���H�}>�`ĂO�����}����@�\� '��@h���p�����Y��|H�#2�Y���~_���	�"��"(�&�r�Y����y��9�J��Ņ��q/3�/�/��������I�F�^���%��gp�! ����#�0��!���/5�����$$$�����8�N#���?7��#E�o���x�j�䂈4�6��N
 �\u<beE�.α��UJe��LM���]�r��\��5�R�\��f+��b�j�ֱ\�2�+]�v8�Z8�8�8�8�8�8�8�8�ŋ,X�b�h�v��gc�b�h�8�N�*T�2eJ�*T�R�ɓ&L�2dɓ&@��I�E

����������(P�B�
@P�AB�`OOOOOOOOOOOQFTTTOOOOQQFFQQQQFFTTO`NOO2==Q1=2
)P�\8$��t>�N�g@1#���~��	��C��I��q��ߠĎ�`bGP����E��t?DA�B7888;��$�}��o���4	�4"&�y<�Bn�3��4l���}���=_���f�	���G��#�����ء�<P�(�l膈H�(N&�Cy�*)����kCCC*J�Jp��f��젿�Y#�WXBgUX@A7@l@oAAB766^^kkooooHH555aaaaaa000q8�\F���"R�����Q"! /$��/6���@�Ý��Ihbd��\�qC�J�pQC�Ru�a��-�je,Gb�j�,X�Z�u�W&L���nݎ:իGq�q�q�q�q�q�q�q�.\�r�˖�wnݻ,�u�V�q��ӥJ�&L�R�J�*T�R�J�*T�2d�)��(�AX�������� @�
((P�	��������	�����*,	��������*�FJ����)��HCCTO
��d�}>�D_o�8;���~��C���t>�Oכ�� �}>�DDD_d��0����"�u	>�o�Б#���t:o����&�{�<���D�@B.��k*��|H��D#7	Dp�)���@�L�f����p")�=dƄ�RP(q54g#3mÂ8��׍LP�͍����ө&�ݬ�UC�E�2fbə��*"�!�;;:**
����������[{{zBBBBBA��	��YD�Aq�, �����g�s�sV@ڪ�cu��͹9�_H�]#o�X	�ɝL.�je,G\�*f)��X�dɗ.\���,X�Z�u�W.\���n�u�V�8�8�8�8�8�8�8�8�\�r�˗-Z8�ݻvY��X�Z8�:T�N�*T�ӧN�:t�R�J�*T�2dɐ (S QB�

���������@� @P�AB�`NNNNNNNN
������(P�X���ѕ�Ӓ�'��

d�Y��q��N�G@8���H&�{	���@��w��03�H��$$�$t<��o7@3��H�u	>����D_��`gC���y�_��bGS��HH�}��O�0��5�H�s[p
#Ĉ`ll�8'���DU��{��![??�̭�Y��s+�,*���4+�4�9���\�*'�������HآH�oų	�p�(-k쨈��������訨HHHF����ck���mmmm���			�y�����qBoo7q#������������3��,+�8�I[��G9"����J,��QQ���&@�T���L�JT˓.bŊիGZ����V�q�Z���q�q�q�q�q�q�q�u˗.\�r�G۷n�;k�Gq�J�)ӧJ�:t�ӧN�*T�R�J�&L�2

Q��
(P�B� @� (P��B�00000000
(QB�
((P�
**)���'���(�FTC )o|Y-��/Fnf�̑��		:�������t:�D�΢GC���$${���O�17И��I�HHHH�t: �O���I�$$�}��@�כ���zg?8.�F?ۇ�6�F"8$}���	��������k8!�i>���c�u'���*G(�(���O+�-+���誦����#�G���op�
 �8H��+*����*���������訨(&������ccck��mmmi�e�f���`�~kkk7kko675H^47H56BA7H67(��XY'WK�tPc���\0�*U�]���\ul��%b;�X�Z�h�bŋ��:իX�b8�8�8�8�8�8�8�8�ŋ,X�b�h�v��gc�b�h�8�R�Jt�ҧN�:t�ӧN�:t�Ӥɓ&@��AE @���B�
(P� @�
(V �B�
(P�B�@�B�
��E9�(P����#�����+��2~\�n��>DHep��\��b"o`7��4�u:�7��;���$y>BOg�! ��E��t����M�$�t<�n0w�3���y��o�@3���hA"����q8�F�Z��0�X�l��r(��ʃY1�ɕ��_���
�9��c�ccB�j�!��҂��҂�J���a���XR�
ņ![��˥��|��p ��Y?d슟��J��M�-��*�����訨((HHHF����ccch�&�Q�S��
�����*[y�:+z��"�Z+
)�A�
�Z*B:����Ϊ��6rx�
��F%O&��2��V�s,V�Z8�b�h㎵j�,X�q�q�q�q�q�q�q�q�Z�jիV�Z�qݻv쳱ֱZ�q�u*R�Jt�ԩR�J�*S�N�:t��dɓ @P���&@PQB�
(P�B�
(P��

+ P�B�
+ P��&(PP�X�
�b\�z,���r�n�q?�-�p�`�[6͔!����������}�� 4	��{(4��� �ϱ'S�E�x���زf�p�9��A��@``b@gC���t:B E++#eŸ�7��P���'<Y8�g�O�E!���i^� �����*cE���9��b)�::�"y��Cz"�!��cca��U�����'�#13&�g>A�>c'��>������ ,�2�������""   3��������!!��3��3������� �3����"�����3���#�"��8�V���Л׍�UW�,�
zz K��t@*x�2a�'�Lus,V�Z;�ֱb�wkV�bŊ�Î8�8�8�8�8�8�8�8�ݻv�۷kV�;�nݖv:�+V�8㎥JT�N�:�*T�R�Jt�ӧN�:L�2d
Qd�

(P�B�
(P�B�
@P�AB�`(P�B�
N``
(�b��
������(�q�pc��U\�o�P��-�rdH����n[����,�4�g-��Ƥf��a"3L������D"�,#l��	Aq7'�� �Sa���cQ�t  i��p�<��G���q8��X\L-hCh��b>|�(�C�I2d���9
0n
)��kkҹ�⼄�C��6��q|\��BWU9@GgA747Zt�ȲV�P-�Y1"�&"��τP'��?d�<�ۭ���쬪�-������������訨((HHF����(��&�(G��f��f��&�h(Cf�,�n!�Fsvq��s�!�F�D�u��stU�tVv�Q�d�g:P�r�*��S@��D��˘�b�j�ݎ����Z�k,W.q�q�q�q�q�q�q�q�,X�bŋZ�qݻv쳱ֱZ�q�u*T�R�J��R�:t�T�N�:T�Rdɓ&L�2
(P�B�
(QB�
(P�B�
(P�	�9<SpRgJ�````NOFT �^ �lo8���	��y�qaa8��'�AD�D#/0����$C��#2��@Sr͂�lۂ�,�,�3,��p�'��}�%6͂٦e�8N,�(J��>϶b� ����ZY�{y�(D(���#f�����EusFl��<O�P"�<�ፉ��1�����%��*���ƀ��n�6l��6l��6xо����ʬ����e<�5g��F�����
,��v}E>N2Yd���(4�94����+������������  #��������!!!�������������"���������3��������������������������2��	D\fclؕ��C\�z��$ +L��UÐ1JT���ұ[�R�p��Ǖ]L��Z�s��v����k�֭vX�gn֮bX���V�Z�J�*T�R�J��R�:u*S�N�*T�2dɓ&L��

P�B�
(P�B�
(P�B�
(P�eJ�&L�T�Db���DQҥ�E,���ST����������`�`8�Yf��|�D"��!E}��D?-�������n[��fٶl�L�4�l�,�3,�2̳L�4����"ٳ��Gے!����CS�!�����lr��q#�ECœ��_�|�;���1��x�0��'�%t�f���AB5|M���[UYh爆������O
�-O���N�k"2�N|`p2�z|0�b��8|";�"�w;����A���ʪ�����r�x��������Ί�������nn�����������n���Ύ�Ί��Ύ����������������hhhhhhhhh�l��z96qG_-�ˀA47S�
�h�e�kW):�u��G*�*�r���,X�J�r�,FV�Z8�Z�h��jգ�,X��r��;q��8�T�R�J�)��R�*T�R�:t�R�ɓ&L�2dɐ @P�B�
(P�D @� @��*T�II�`L��� �� �t���׆��ח���׍͍X[��M[���LMM�����D�Q8�טW՚�%��~(�H�b!>
|_��~_��n��n�fٶ�n[���~_���~[���-��D"2N&A�ٲ�X�
*���r�'��,�d铠�>c�a�Fs����,]�5?�Y��QRG7F[PY)_ihA?�=9",�/����"�$5�,������E�d珉E��S,.h��Ɉ�����J�~<⛗��֧8ћ+j��B��+*�Kaʺ��"���::;;:**











�:*

*)�!�;;;:;;;;;;;;9���������"�b�:A���%`�s�О�0_C&�OwF%[L�ab��o6J�
V�=Qv��˖��b;����Z�q�v+��X�떎��ŝ�֭Z;��u*T�R�J�ɔ�R�*T�N�:T�Rdɓ&L�2�ɓ @� @� @�dɓ&L�2dɐ
���A�==�P����S.I4k056g@AAB76^GE7kk^ok^^oHkA5q8�E�z	��I���d2��� �q(���b1���@�S���/����/�|>��b0|�Q0aq7���͐PW�O��_.�v䊇���~��NϬ�S�fU]@��v��ؤ��A��8��P��!�B�@������opN��(�H����o��k?�'1�i���Tʌ�8s���1���d�'N}v3#��!���eg����Ֆ��VUT�Õu���DDDDttvvvvvvvvvvvvuu�CFtTTS��DtvttttttttttDDDDDDDFut�D$#tSDw;t�a�z��xT.y�1ED��U�  �P�{���r�b��vzh��f+]�,�u���b�c��GvXab�ݖv�s�GqԩR�J�*T�R�*T�R�:t�R�J�*T�R�J�*T�2d	�&L�2dɓ&L�2dɓ&L�2d�
 @�����D�%:�̰��Ί��΂��Ί��nll�h�n��nl6ll6��l�΄����ސ�oHgjI5q�F,,,.'���8�J'����F#��b1�F#����D�Q8�N.&C� ��Q5a7^k7ABgG4XmVhGfY����d�%ߋ~��RG��#�ȲgY��5vA|���d�K��&d��r�䊜�R<EH�2|'��܂���p��|��8�' �!��QT<�,������ԧ �Q'��Gc�H���,�d��3�nN��g'����Ֆ��UT�Õuu������DDCCCDtttttttt���vvvs�s�DttsCCCCCCCDDDDDDDDDDDDDDDDD�ttDU�Fq�VA��5��66ie=��¦����f��<1�m�uJ�0gqrr��G�k��� �2�,GvY��ݖ,�tŮ�,���:�*T�R�JT�R�:T�T�N�*T�R�J�*T�ӧJ�*L�R�J�*T�2dɓ&L� @�zpReN�:�*�˒�Q&b�s�"��"  3������������ �������������"����/7�3�+"2�R����RMXLN'���d2'�!��?��N'���q�0������YЍ���UQ�G��,�~#'��(�)���m� H�1�h��'�x��Y�&C ݐ0�`sc$Q��� ����$3�+6 66 ����B�����R�DfK$c��S�X?�6�}��yI@Á8N�8H0�ӝ�f������ڲоʪ���rr�����xxx�������������ذ�hh����x�hh��������������������������hh��hr���Ί��lj�؊��������n�+0�+FBy0��VYL�ZW��Ԏu\����L1���*�֝F{��J��똭q֭R28�e�V�R�J�*T�:t�R�I�J��ӥJ�*T�R�J�J��ӥJ�*T�R�J�&L�2dɓ(P�B�
N``
������Ry����Y4BE<IG4DD@@<X@@DDD<<<V9EGDGg444GEAg<lD4EEggA7BlYUXE6E67BAB6^o^^koHHH555aaa00aa5HHooHoookkk^ok^BGDDAD9XWemYi3m^nN��,ˁ4�L�?�w ��Bd�FȈMl��iV�ۈ�jސj���"�ݡ7�#����Y�a�[r��nnhx����r��6�Q}&�����%#*Z��H���7�o�E��Q@?	���M��k��)PrzxjiiYh_eeIIIlll99WWWXX<<<DDDDDDDDl9XD@@@@<D@44@D<@@@@@@@@DDDDDDDD@@@@@@@@4GA7gXDA6D@GD4G<GkEXgAg7kA5WiEAAEI	I^mjUADE<GBGU|�?� ����_*��wI4�����5�Ř
&uJe�V�b���B�wZŋ*T�R�J�%J�*L�	R�:t�R�N�:t�өR�:t�R�J�*T�R�ɓ&L�2b�
(P�D�0#����b2GKJ�*:"º����JJ�:9��¹�bJIKb*��:��!�:���:9��:
	�J��x�m����y���lmyyy�����!!!��xllll������	�a\��%%����`�����A>����	��>���� �F,u��
a0A6gJ�������j����8I��8Ts���ZC6ͯ0��l�nn��Ԡ����h΀:b0��h�#����"7��!��DN'�>�p�O��p'��<�En��՜���[VZ�UUURR[NU���U�PMАV��Y��OM�Б����VN[_(H-�
��(��(�)),&��-f�	�*��eS�^J�������	T�\Ŋ���%=:1j�˗)R�J�*T�J��ӥJ�:t�ӧN�:t�ӧN�J��ӥJ�R�*T�N�*(�d�)*9�(V	N�8�Y[NNNNNNNNNNNNNNNRV�[J[NP[N[����P�O�QPPPPPPPPP�����͍������А���M��U�^�]!�œ̗d�����l<� ���~^�� hۡ � ټ�m!ƹ1ף#e䃊AɊP�R#�i�)�D3lĎe�4p��|���)ViU4V
����:QJ,��]	a� �DM�q>�g�|
}9��d��%Ϥ8L�cE/"��3�kk�R�ʪ��JJKccca��ʺ��""""""""��""º��������c��C;a�********


**+;:*+;;::::::::::::���#:)�a�:�J�º"""""""":::::::;:;:	�ȁ3�G*�� �yu0E�e,R���	_W
:Y��*T�R�J��R�:t�S�N�:t�ӧN�:t�ԩR�:t�U*R�:t�Ҥɕ:T*y���QI������M)')))))))))))))))),��������	*��.uUUUUUUUV�UUuu����V��E�u�w�5SCńuuu��CCDvvvvvvvvvtTTT$$$TTTtTtEs�$TE���TG�0e Q8� �'��N��~0�nM
^�`��H&�f��F�o�#�����9�2���Y1r�s��>Ϳ%1�|H�Q�չpXP���AD`P-�?����J!��Oe�Z�Q�
�9�!��	\���>~Y#$>!�2�. >�K���!����ixzxmhe_UUUUIIll9999WWWXDDDDDDDDWXD44DXW@@@@@@@@44444444GGGGGGGG4gUm@A4EEEEEEEEEAAAEEEggEEEggGGGGGGGGGGGE7BG4gGDE44gEgGg@@@@@@@@GGGGGGGGEgE4GAP%L �Y@gg^gg �'8�J��X�dx�U?��]�bd �J�*T�R�*T�N�*�*T�R�Jt�ӧN�:�)ӧJ�*�)ӧJ�*t�P��N`OF1n��(9,����������������������������������9��VUYZ���YW�NU�\��Y[�[U�����NOUT�NQ_"N�B���d�����@�p y2y���6z�u'XG�$��Sft��A��h�#e�ǝ�؋8*.���"��w�C�d���(d��|)d�����#�YA>,��%��H��FL�L�+�$��_�&��rhx��n�&"�6�G�Mϝ�9���(,����8����Yᵡ�}}UUU%%%���]]]aa`���������`� �� �`���������������ѝ��������!A���	�����!����aa�����������)؊*(������h�4,�)PM ����*��7���*T�R�J�)R�:t�T�R�J�)ӧN�:t�S�N�*T�ӥJ�&L��
*��%Qu:U�URW�[VVZ��[[[[[[[[[[[[[[[Z������������ZZZZZZZZZZ�ZU��[W�W�Nf�VS����VUUT����������Ó��uu����Ņ�uuutu�V����&�VV�M$��n >	�#���?�,�g� ����	UU��T��X��9���,�Ԟ��b��R���6�2���!��
!���	��!��y��j�� �˓`�톇���,�j�u��L�fY�O1���)���,�wۄ͕�����%%%�����aaa`��a��a��������ф��Am�		����y����my�������������������m	��u�y�����y		���DB764_ ���o�T�R�J�*T�R�)өR�J�*T�N�:t�ӧN�*T�2dɓ&@��D�00
���rmmjzjxxxxxV3jjjjjjjjxxxxxxxxxxxxxxxxxxjjxVVrxxxxxxxxjxiYjPViimjzi_zhehU_rYYYYhhhh________eeeUUUIIlIIIUUUelIee_hixe)|�g�('�|'��������"p#�D`���s���C�u�C�T ��X�
w��v$�n�5��)�XQ�H'�%LLQV)��b�s�S&%/�F{��JURɤ���� ��lh>��"�Ď�?d��A�"*���y��e��}}T����]]]\���� ѝ�� 񝝝������y	U�%�				�����������ݝ��f׏���QQQQQQQY��������F��ז@CW�PM�����Y�QY�F��)���/�*���-g�*T�R�J�ɔ�R�*U*T�R�J��N�:t�ӧJ�&L�2
((T�iJ�?�ne�֗���'���������������''''''''���������'���5�''''''''���ע�e����g��� pj�kk��KKKKKKKKkkkkkkkj���CCB������CB�˙A���A��n��Ȱ�P�Q@?����8�|@� }��':ehff$���U�D�S�tF����WHn����m�7 \�~��?�B�#N'��3���{����YI�ڜƸ�+�Y�,Q��:+;z;Q�YU��͇���>k�s�(@��6|Ÿ���%��aaa`�� �����������								����m							��				����������������� "����������������#�� �"��#������������!��"�$7���0��$�)R�J�*T�L�J��R�R�J�*T�:t�ӧN�*T�2d
(PP�	�*�!��w'�����և����''��'''''''%eeeeeeeeeeeeeeeg#5g�f�Kk�����������Q�t�eA��Y��4%�Ҳ�ff���������������������ڲ��������Ҳʾ��)ia>'�>a�#�>�1����� �p��  � R1��D?��#���������"�4 ���eBI>�uEA�;{�J�29pC��@���<�K,�>|P3'O��\<� �O�G�	A#��n[�U�.�B]�,�"Hrٰ, !��5��,4 2�����662�� ���-�����������������������訬�((((((((HHHHHHHH(((((((&�KƆ���HHHHHHHF���HH(((HH(((����������������(&��興�������������������&��HJ������&���h,�m�kȇ�ml��k���HK��f���T�R�J�)�&R�JT�T�R�J�'N�:t�ӥJ�&L��
�����I �j���KKÓ��S�ћ��R��������䠠������ffffffff��3z3s4�+++++++��99Ɯ�m-�OOB%�w&֕�Y���������������ᩩ������e���������A��f 0���O���t}N�w���h��H&� r6�xxڰ�ʾ�����xrxЂ2J�UpNԭ�ҳ�҅h#�ɒ�Ǐ�Gҟ���_�__'���R~>	�?��'O����ـ_��u��E�;v.�ND^G^6^qZIGµ��*Mo�c��� ����  #��� #������������3���� !!!!!!!!!!!!!!!! ���������/5����!!!!!!!!���!! ��! ���������������!3���"��*�$"� ������������������3����3��� !3�!3�� �� #���3�5����\�2e*T�\�2e*T�L�2�)R�R�*S�N�*(+ QD��*(�'��<�*�J�O
��������














fffffffe%%%%%%%.g9������Ü!���A�AY��jzt�=8A����ޝ#NMJoMNJ�NNNNNNNNJ��NOOOOOOOOOFov���������@<���Y���>k�L��J��� ��Y��CkCB��C*�J��";J��WH}�^/E���{�3�H�07�������ϯ>��^>�}5��0C�w����~0} y߁p�L������늦Ju8���
��{4n?/��:䣼/!��F`L��b�)���M�PM������QY��������QQQQQQQMPQQM��PPPPPPPP����PPQQ��Z��P�QQQQQQQQPP����QP���Ѝ͍͐�Y���������QY��������������������QQQQQQQQQY������������������������PPPPPPPY�QQPPPP�����.\�2�*W.L�J�*S&R�JT�R�:t�R�SӅ 9E=9�*y���rxPs��++++++++��������������������������w;���s���%&e%.ue�5b�1�ә��s�(:@��g����3rVp��^��U���������������������������D�
{�� ns2�f׆����3�LXĚ���c�㓖�ֆ����UT�Utv�`q�GE>(�笃���T�����Y��";��L�ߎO�� �L~d�Gy��%�JO�/�!������K��@�,�|"*&���殊��
�6d8�P�G�A|�q�%���HT�\MQ��0J���9��;;;;:***+;;;;;;;:********:J
*	��










**�*��;:*******+:*

+9��9�
�:	�:;9�:::::::;;;::9��������������:;;;;;;;;;;;::::::::;;;;;;;;:::::::::::::::::;;;:***;;::�˓&R�Jdɓ)R�*�*R�:t�R�I� @�2{ P�	�)���!�7	K�KK���R�ffffffffRRRRRRRR�s9��g3���s9��g3���s9��g3���s9��g3���)rVn�7F�/'�3u�Y��}�����!�"��7;��AX̥AAAAAAA@��AAAYYYAYYY����Aΰ�[,�|r�R��D��˿�6/6�,��44/����"���]�Rf��6�����Fl�7~)�3�Oǳ�ǄwY�_�ߌߌߎ���^#�}5��%3�gי)3(�⏘v`�}J�� 0����U8�R��Qd������k'N'�Y(�԰bd����n�nh�������������������������؄��n�������������������n�؊n�h���������Ί���Ύh�������hhhh��h�hhhhhhhh�hhh����������������hhh�hhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhh��������hhh������Ύ��r�ɔ�R�2e*R�J�)ӧJ�*@�B�
(*rz��zr�p�h�YAYA��|������������w;���s�_/�����|�_/�����|�_/�����|�[���������s9�!ד�����44�}:�bmґ�IIHә��|���%%%%%%%%%&ffj

j


����
.��œ:��b�A��������W�YW�W���U[OВXA�,dhRu�ܿ �m�Q��O�����07��߂3�K~
Gx�a����O��_~<||?ϥ�K~8d��<`��/ƈ�d���03��8��จ��^�i��>8AN#!d�j�L��!�	J����tt$sD$$TTTTTTTTTTTTTTTTVv�$TT#�TTTTTTTTTTTVvvvtu�Tt#DTTTTTTTTDtttsDFt��DCE�sE�DDtDC����������������DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC���������DDDCCCCE˗&L�J��T�J�)ӧJ�&L�1B�
���@�Iʅ�����Y@���n����뜥��s9��g3���n�[���t               !��|�_/�����t�]#A�7�@C�K���s�?�Z��/�� ;� ��i��rPp�9��g%f���s���w9III����������������J�  U��1L�(�̋�؃X��,uP]x�]%U%UUU%�]`�����\�=}����Q|^"�ψ-A���>�����'̟����������_���)?�~
}0��0W�'��ƙ(d����(��ȱG\��	�8�V�8��0-�(���i{'J�R.~��,U<Y4��Y�����		�����������%�����$� ���%�\�� ��U\������������aaa]]]]]]]]]]]]]]]]aa`�]]]]]]]]aaaaaaaaaaaaaaaaaaaaaaa`��������]]]a`���r�ɓ)R�J�)R�:t�2d� (PP�X�X	�Ou9��\�r�9I��K��4�n�[���u�4444444444444444�n�<��N��;���U<s�4���F�]/�����y4(���9��\�Ng��3���s���w9III��������������J�K�k`BQ�;ZXc�+y�ڗv3�ᇍ��*�'''*������!��@� ~#8-�����|�G���?�P�<EO�����E% �J�K� |�U�_���LE�l�\� ť�7!��,�\=����Ÿ4��:L���0�#L�����l�n6n���n����Ύ��������Ύ�������h��hh�ʈ�������������xxx�lή�hx�����������xxxx���ΰ�خ�xr����r��rrrrrrrr��rr����������������rr����������rrrrrrrrrrrrrrrr�������������������rrr�������r�ɔ�R�JT�N�:L��
((P�	�����1�9K��44�s����g;��444444444�t�].�K��44444444�|�_/����R�y8@�!w�t ���HE�I��t?�`o�8Ӆ��s+(�9�[\�%%%%%%%&ffj


��


��NNL�/�!�2˙޴�R���(��#�R�M*\��x�xxx���x�h���hnxQ};,)��̇�O�X|=G�A��y��>vJ������b�Dt�/��$y�Cœ�' 2y����)(/��_	�Y�pH��ZJ�����nY�m�i1\T�3�S�������X�s���!�!! ����         2��" ,��,,,+�����!,�������������,+�������*���2�RRVVRRRRRRR[RRUURRRRRRRRUURRR[UUUUUUURRRRRRRR[NNNNNNN[UURR[.\�2�*T�J�)ӧH (P��E

+T��3�!��s7F�#A�'�C���t�].�K���|�_/�����3s�<� N���';���Is�����`�!�� K�Ҭ�}>ZU���B��.v�����������35eeeeeg'''�;�JJ��å���eT������䒥t����CTCDDDDDDCDvtTt#��Ы,��8�'��pO4����p�d����	#�Ġ��p�|�pC��d〔������Y (������O�pͳojB��,��fߐ[�Ԇ���L���R��h`:��r�Z�+:

:9�"""""""""����#i��������º����cccj)�!��B�JJJJJJJKcaʺ��cb���cCi���yeUU�]��������%%%%UUU�UUUUUUUU�UUU%%%%��������UUUUUUUU%%%%%%%%��������UUUUUUUU���UU%%%%%UUrdɔ�R��Rdɐ @����Υ&��+p���44�3|�_j�N`��˒������y>] Ng������� �u�H�Pn��� ���� BGC�� ����\b̨�u�HC��n������������(((����+(+<4�6��2��,�P�	�79���BJ;���#-:,�6^AUE@gg@X@76A5m|L��c��(O��������xX�!�OnCœ��d����Nd��3,Ӏ����8�a^E@Edg��J ��� Ud�|H�f�q���S18śnJ�R�`
������'�J�lnn����Ύ�hhh���x�����������������rr�ʪ�ʪ��r�ؒ�������ʾ�������ʾ�����ڰԾְ�6���Ԫ���nΰ���ڲ���������������������������������������о������������������������������ʾ����ʪ������J�)R�:T�2d ���(�2d*TR����n�\ N�����������������������������������y9��N�3�!��z3y+?]Nr������}�C\�E @OK @N��C���}����`)-җ��@@@@C���)))))))))3PPPP3)hmzVPVxjPjx)r_r�R��s����xr��؀�v1���N� ����! 3�� #��!5�ߖJ,iȤY�F(���;�J��p�d�������|,�����O����|��8�Y��X���v���?�����ec����4�dtꐤ�C��!�¬AE΄����Ύ�������xx����rr��rrrrrrrrھ����о�о��ʾ�����������������в��������UDzEHXA9rm_jme_hmjxzziiiiiiiiiiiiiiiiiiiiiiiiYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYhhhhhhhhhhhhhhhhYYYhh___mmmmJ�)ӥJ�&L�2
 @�X�
`Q=y>J\ΐ��hhhhhhhhhhhhhhhhhhhhhhhhhhhh !��s�BN��u��s�4<9���7���)Up���!�`��b������f�9,:]%+� Ng'8�I���n�:F��w;������������A@̤����YAY�A���e�	���ǃf��+*����c�\����`g4GG4D@GE7lg~)��L]���D��(��f�]����*�'�"�%��Y�߁d���Œ�Ň�<,�(�88P�>EN �CĠ���|��3A���jZ������ə��P�#&LęU�색���Y����!�;:9��"!���º���ccbJJ���++++++++�J��KSSkSSKkkKKSKKKKKKKK��������KKKSSSSR���%��~gEePzjzj3PzjjxrVrrrrrrrrrrrrrrrrxxxxxxxxiiiiiiiijjjjjjjjiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiijjiimmmmiiii:T�Rdɐ&L��
JT�VDʰ���@o ���@����s�>_% cNa12�� ͩ}U�Y��|���	���'k����|�<�O'BK���zx{,��J\�o�a� 0!�7˘!�4�))s9��w;���s��L��\�NJ���OMO
�M�M�'S�� 񕱡��$�%���c���1B(�/+� , #��������aS�Fe�q8���my��4϶�E��<P���fO�!E��j���l��qnN,�nH��l��@pH̃�r���p;�D ��J���v�s�S�0������ ����",+���66$����������44,��������<6��=<5=<<55<=9========++++++++99=<554����ZV��T�ܕU���������������������������������������������������������������&L�	� @P�ASӂ� L���L!��t�������-ґ����������������������������������n�[�g&��V���u�	��)t�?@ۮ� '���!��}��8�!��ﰗ�K�hD@�M��s�ۡ�3���s���w;���)3333)s�++++99=54�<56�95*�"64,��54*�������b1rӨn�f�v�DU��SC�r(>D=O�,��̲'C���:b��pY zEO���#��|�	BP��-�fH���$T������8���?6��,�����z��4�#̐=~B�\Ě�%���H���(��g'-�)*�������+-���---/
�M-/OOOOJ�
��������






j
OOME.@�
��O�	K�A�������f��Ԡ�����������������������������������������������������������������������������������T�2d @�B�
��4�W�0���|�:@��O'H����������������������������@C��x��s�:_J.M
��'�n3���_x{������N�K���n�� 8D]A���#0"�;���@hB�I��� i��s9��g3���s��L��\�s5eg''&��������'����T��T��V��U�S��F.Zt$E��6AXl<Bg9WAd���BQ q��Q�n#�Ő`Q"!/����̀��?,���n�Dd��gď�b,�d�y�_�_��	�8 �������r�q�(�ϰ����E-:.ބ�����Ί���r�ʾ�в��������������������������f���䠬��������fffffffffffffffff�))3PVVr3hn�ߣK�'#Of�Ҫ�kћt!�R�����������������RRRRRRRRffffffffffffffffffffffffffffffffffffffffffffffffRRfff�������T�Rd� @��B��
@*�����A��|�<�Af��hhi��|�UZ�DJTo�g9KR��X�� H�����(=�������|�W�A��I[���3Л�ЛÝ��R��f�y9��g3���s9��r�32�;��R���䬬�������ڮ�f�����lIemji_lu;�b�D �͑URNQ��UJ.G|��2Ij�N@pMX\N#��`w[��p y?������"�:~#�����߅��2y���FbG������� �g��(\���2�k2�H�~���� ES\�i0�vtu�sÓ��V�Օ��֖����������'''%eee�J��K��R����f�s����������w;���s���w;��������$y<=+9���w�7;u��s9�JJJJJJJJJJJJJJJ\�w;���s���w;���s����������JJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJ\�%%&fffj


J�*L�
((P���7�C�h	��t�>B��.g0C�hhhhhhhhhhhhhhhhhhhhhhhhhhhh !��)~Z��^a
ϗ˒ʪE|4	��s<���-�8h����t�<�O��P8���_A�-��N�'&�6����� !���s9��g3���))))s���&j�NJ���jJ�*�.fՃ������&�����S��F.Zt$�M�Qxl<GlPlf`�Y��X4�7F`X~Z�M\L+�B��@O��.|���88$p��,�-�HAkPO��f�#1d�Y�#��B缜K��g�1��$XnO�jV�0r��tsEusŖ���ev֖���������'%eeeeee335 ����|�[�


.v�䤤��������n�[���u��s9����t	��rmt��:Z�����&뜥A@���s9��g3���s9��g3���s9��g3���s9��g3���33333333))))))))))))))))))))))))))))))))s��JJL���	�&L�����E��'H�@@@�@@@@@@@@@@@@@@@C���t�].�H@@@@@@@@���������������ӅT���t�\��';tͥ��E�R�q���/�Hh3����y=����m�/5c򖀇�uά��Vt��\�Ó��p�<(7F��w;���������������ɥ�R�в�����Ҳ����-;J� ޮҎt��	�����> �0f�� 9�"CY�ٺA�X t�8$[�H��>���� �@(�q?���3����P�G�fJ�����XOP���ߔG�:�3 ��&�b�G<@eeYmmmiijjjzzzrrrVVVVVVPP33s���w;���s9��r��37J��u��)ghs>\�g3�!��)mYr|�������J�ɺ�n���e`��˙�4�}=9�Z���ϗ����|�_/�����|�_/�����|�_/��u��s9����u��n�[���u��n�[���u��n�[���u��n�[�g3���s9��g3���s9����u��n�[�w;��T�D	�R��^�q��#@O!����                  hhhhhhhh        hhhhhhhhhhhhhhhh!��֪�n��M�H��H����t9���@L��� ��k���m�s8�-mg1"��u����rlIriV3U3s462���F��g3���s�����+++++++6�<<((++9�V^�Z��ŧd���Ư�e�LP;fE�Dnes�x�`U�A���X)e���^��� �XzP�/�$"��EH�pl�q0�/5�[�!��np�e�\��A����� ����
U"���
&�*�#�42�/�����55<<9999+++(+(((������w;���s���g3���s��_.�3�AT�� i��|�B���Fe/
'�C��!��|�Lۡ�H@@@�K�I�Xͺ�|�_/����444�|�_/�����|�_/�����|�_/�����|�_/�����|�[���u��n�\�g3���s9����u��n�\�g3��ӥE'�����O�9��h!��|�B����������������.�K���t�].�K���t�\�s��8iI�����R�y�Ą�\�$�`$s�A���b��#��I+��h��}��P rDIV)u9�B��Ї��̒��Ҡ�t�>[���u��s9��s33333330�5g3uY��驩�Y���b0bX��!K"��ID�Nh]�R�nފ����Y�QO�����JA�R<G�>GpH�>'�
)�6����\N	�#��'������LɊ�l�$��2U����� � T�T�S�Ulm_YjjxxzzzzVVVPP333333))s���g3���s9��g3u��|�B-Ѡ&�K���t	��t�\ϑ���:������5��f�y:_.a��K��44�9Xn��#CCCCCCCCCCCCCCCA'����t�>_/�����|�_/�����|�_/�����|�[���T�J� ����-�����4�n�[���������������������������K���t�].�K���t�].�K���t�].�����R�)IgUVzt���
��5�3k��F)=zp� �@�!��7�"3K�h��5��Y�$�Pt��(<��_&jo�����y>_/��u��s���w;���s�\�M�
k-E&nE��� �����	K�m�;�� �lo6BD$�ޑ��[Y�ۢ&E��pH�d̐�8�8~8�3g�>����p2*GωA#��E_��8	@"2�A��a��y	��u:Ŗ��r�֒ �$�9==999+++�������w;���s9�������|�_/����44�t�L�ΐ�����k��4�y:F�/'��R�t����Ӥhh4	��y8C@�^�_! o'����y<�N�K���t�].�K���t�] @O'����t�0'���U��!��C���n�[��������������������������������y<�O'����y<�O'����y<�O!ș�s�!�H�Wk4mn��@��2�t��f��_rxhm ����YDD��CK/���+�$E��s=��ᮠ�F�G����s9� bnH����t��.��������u��n�[��;�HC��u��R�r������Z@���n��	0D���W�Q��eu�ՔD%��H`��3%&f!�-��\,��~3,�D�m�
0#����
pAEUqg	�uU] �m3*�{H3��$��r�֒ �$��++(((�����w3���n�[�����44444444444�t�^@ng0@@k�	��|�^COg�44	e�A�4�y>\#An;�5��|���A��                '����y<�O'����t�<�O'����y<�O'����y<�O'����y<�O'����y:].�K���t�].�K���t�].�K���t��:B!������ hh!��|�B�.�K���t�].�K���t�].�K���t�]/'����y<�@@@@@@@@@@@@@@@@BA BA� Į�2�u��IX	y/�]e���es�2�$Rʪ�� �I@��z�ap�� _cO��4`���H@��I��)~��+O��h	��t�� @O'����t�>T/���+�βrhj��&u��y�����˅���^�U�I%��NR[M�-�Ĩ��h��Fe�fٰ[6p�&�Ő�`�jD(�[�-�2c�Ɏ	��R�PO������5d�'K�ɣtq���Z��/�K�斕2U+_ʩ//fe%%.w;���n�_!CCN�K���t�].�K���t�F���K� ��p�F���CC\!�oa1�&����n��#N�����{>�n��E��0h���hhhhhhhk���p�\.���t�]#CN���p�\.���p�\.���p�\.���p�\ @@@@@@@O'����y<�O'����y<�O'���H"�s9� Ob�3�i��y<�/�������t�].�K���t�].�K���y<�O'����p�\.���p�\.�K�� �Ct��b�j�!�@���D��h�� �}���:����A��J����z�pC@h���k��4&�n�/�9�M�����{=�@�N7���y=�O����"8�J��ij']�,��X]<(q Л���#��46/���V\�
	@��U@љ\ ��C��ل�������o��f_��"ٶ��8[� |����>ܜ_�bG�	�#�3��a�1i׆ƅ�W!��T��V�,�94�9��w;���n�B������.�K���y<�O'����p�<��-���4	��y��C^��NgK�L4	��gHYz)n�_A�O1'��h��i�B��4�@44444445��p�\.�5��p���������������������������������\.���p�\.���p�:^@O'H�Ӥ	��|���� NK���t�].�K���t�].�               '���p�\.���p�\.�P�p 2� �������{�8U	�/��wXk٩]���zO,��}���p�����G6YX~����"�N��4��^Bb"``O'hhk���t�].�K��f�s9���b&,�s:�T�/�pũĮ�W�0�rK'ne�$�$U�Ƨ������|�v �eDR-�pO�,�!��JZ+c��J
"!��8(�Y#�Df�	Ad�|�|_ �ڒ��&Rؒ����y>�AjFL�]a��Y��s9����t  hhi��t�].�����|��﷓�L��y8^�g���M���}�F���A��K�L��t	��:��@��71����{=��g����p�\.���p�\.���p�\/'����y<�O'����y<�O'����y<�@@@@@@@@N���p�\!��������```````og����{=���'�Mξ��u?�	 ɺ�.P�̀ ���49%~���������&d�EޖD����H4�.� ��1v�08hC���8\���L�%Y��|��:��	*�g����p�\ @@O'�t !��}��>[�%F-vUk����	�O8k����XhUmrl�\�f�̸����J,�ɟ��8_�� �o�Px���2G��/�p �(�����>��p7f�E�n�$y���Z�@��t�9�j��`8��mjӣ<��Z��[��g9����t�].���h��t��!�o`01'���ڒ�$$p��	��\!�o�3�M��t�(</��<� Ϧ�#���}��	9� �o��袒&&&&&&&&&&&&&&&&&�}���D���������g����{=��g����{=��g����{=���������������������������������CCC@��������������������������������CCCCCCCCCCCCCCC^�g����{=��g����{=�b n��c7���"� ~�������o�p30b��I��q���[F�H?�O@�ngכP3�H!�ō��rUPzDaz?3
8z��44�u	�=:IFo����p��\.    'ɺ�y�ܜ�(i��G*8�@]&IV�.QR��|5��%%U������4��Dp��Be\̡�5ssa�������dٓ�"7-È�q?�׍A`�d��N$C�ѥW��ŌޛYZV\�c7���GR�q�Õg����|�<�.���4	��}<���L��!1!!7��5�"$�p���ϵf�ڳ�S(��5��t	��ۡ�mi�%��t��H&&&&&&&&&&&&&&&&"�}����������������������������������������������g����{��������������������\.���p�\.���p�\.���p�������������������������������������������ANp0g؈0c�LI��$ t�^�78������f ��U�U�J���Hb�ʾ�q����f*�1����[S��̐�y���D��``cOJ�K��H���445��p����� b"i% 鋓إ-[:� ��`��p��S����e��:��(pG@/p�����>|��H���,��\����>��n�FJ�2͸!��~�>$[1|LP_��H��>ٖO0��"�(sS��IJ�(���3�.ؕ\$�Բ�R���y9��`     '���p�	����؈��LE�"���}��@�ϱ��HHI�&�{=��J �'2����{��" .��I�{`��H�Y���xkt�>�o�����}��o�����}���O�1Ј��������������������������������������������������{=��g����{=��g�hhhhhhhhhhhhhhhhhhhhhhhh���{=��g���������������������������H�u	>����/`�G[�I��{>ĀIB�7�s��r�u�Ɠ��2� ����̀Y��q�_*�[c���zr)	1$iY{8�#O��Cu�H�rt����bbb/g�hhhk��"�)zt� &�d,J�Ik��E����x��`=`.3s=2���:��7U_ �($X%QT�/�6E�n	�F78����'�scSFU�S�FtS�V�v�@)�f٦m�#��qp�]C)�NJ^!��d�,�h�#t����%�f����${<��b"og���I��{�9�@Bog��E¬H�t	�9��o�0rA7����R  �y���N�2�a�P�c�  h$��M��}>�O�����}>�O����"�}��ğO�����}>�o�����}��o�����}��o�����}��DDDDDDDDDDDDDDDD�����������������g����{=��g����{=��g����{=��g��LLLLLLLLDDDDDDDE��}��o�����}��o�����}>�O����"�$~�@Πgө��t�:Og�t5��}>Ą�g�ā�!)� ���(��t8_��O1���W���򀬮h J|�ӗ��D�о4&�}����O���LM��{�����!�`�4�G����1pJ����J�(�ӌ�)(l(�v�J��M!���	K��Z��-f��#r�$d̑���8�8a>Dx������B)|��'��C��8�����TeYVF���Jm�7e�B�7��q�����3ep�:@�^�bog���	��y>����_bD��!'ۨL4�&"&�t��^Bn�gS��&�u>���j��O�P��H"&�_emu:�n�:��!�ξ�}:�N�S���u:�N�S���u>���bb/�A!!!!!!!'����}>�O�����}>�O�����}>�O�����}>�O�����}��o�����}��o�����}>�O�����}>�O�!!!!!!!! א�!! 01#�M� ,&H�q�	=�oN�ׁ'�   ��\Hdd�I}�	���$0bA�0C%��1���Q2G�ћ��"�����9�n��H���&�u:�O�А��������p�:DăL��`MM�H ���M� $8�8���xl�"�Yˀ% ШJ�sO�$"�:p7�f�"���H��8�|�p%�2Fl�(N��"_m�pY���/��⼮�pY*G�\e��栁��9KS����f)F�^ ��/'������"�}�������_`bo�'S���}�����#���$y<��:�Ď������7EP}?CU��o���D���&� u�:�															N�'ؘ����u:�N�S��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$�}>�O�����}>�O�����}>�O�����}��o�����}��o�����}��o�����}��o�����}��bBBBBBBBBBBBBBBBBBBBBBBBN�S���u:�D�'����u>[D��@��gK�D��J� y��n��@c%)������iq)a*����<\$�Hr��{�ŋ�owZ��kɵU���3"+<��ϧ����}>�N���DDDLLLLL5�"�t��l�D��Tp��lI�>�	[Ry��HЋ�Is�ɤ45�Q~����P�X�֒D5�����P��f��1�E�m�(Y�Y�͸ �m�fϳ����L�J	�qlf'�"#ޜ�Ԡf�mxbY�e�W:D�\&nuW�Ȉ@���$�}��8��/�1�#�I��{���	O�GS���y9��"@�ĂO�72H���4�UY$~���ۯ`q�����y�	<� DM�_n�```````````````bBGS�LE��$$$$$$$$u:�N�S���u:�N�S���u:�N�S���$$$$$$$$}>�O�����}>�O�����}>�O�����}��o�����}��o�����}��o�����}>�O�!!!!!!!'S���u:�N�!!!!!!!'S���u:�N��C���|��O��  ����H�u���B���g��\1�n�9�=�����I���=�o@1t�AP�0;�}@E��s�Z^
^@�*�D��ȋ�I�$�}��O����""&&$H"�s����b�NB`�c�&�$h�F�7\i��J_g-�g띡����9�O.u�х���d���ɏ�<O�������_��G�p">�H����% P pɓ#�O8���Y�������J���"�9|�>�1RY��a�&�y		�:�F�F��ϧP��E��WP}��ĉ`��u��}>�N�7����4�u?_��GP`i��ar�&$ �y�ބAN����L��$ k}	�:�C���t:�C���t:�bb$�2BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA!!!!!!!!!!!!!!!!!!!!!!!'����u:�N�S���u:�N�S���$$$$$$$$$$$$$$$$u:�N�S���u:��ߡ�w�wؓ�":ȓ��$�t:�`�p!w���"#�5� ֎�%$t �/b�FF{���(��:��Ng8b9H#���t�>�Є�oO���ɛ�E@5�H� p��BBBO���5��$}�����3Ԯֱ`�'OS��������Š�Z�庒 (��X��){�@��nE�!��#�p���<�R)8�#�x��	�8�A�>	�f,�>w�>O�=>N}G����G��rR�lۤF��;�B;h������@0C����H��}��O�А��#�D��XHI�$$&H���y�9���BG;��4�"�y���XP��D^���a��w�Ku��}�<��7�#���y�	�I_������~�_������~�A���������C���t:�C���t:�@01!! 00000001!!!!!!!!!!!!!!! 00000000���H�u:�N�S���u:�N�S��HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH�$$u=�o�J��"�hUu	:C��7����~���!��;�� ���zz��J�,��Y Q\��}0 ��*�g;������Ys:�M���-O�X8����s*�^`ΧS��$$�}8�����'3����q���%Z�p�-J.zbH 1P�7��A��f�{< (�Rb�rq���@PN �L�>�'���O2p�Pd�@�|��X���d������ ����0�����Ϡ����8�>��#�	ɣ6Ys:Pƚ��O7C�lh����7���|�_bo#5W���$$$�u��M�� 78k���&�u��@O�&�"P73���}��@Ѝ��F�of�w	!�H8��40A��<����s�I�� q�>�������~�_������~�_��C���t:�C���t:�C���t:�C��H�t:�C��HHHHHHHHH�$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$t:�C���t:�C���y�B_��B�)�S� ��$ >�OB ���7Az����T���u�����ֱ9{�:�^O4iQd7[��&&�u��Q��].7ؘp���1�R�t	��Υ�'H1!!#���$}�����-B/��Ȱ��ɗ0`낅FFOCO,\J�	u�>���/O繑)��(�c��^�fH��J���_�\	�����*�'œ8������4�5?���D#� �#��ݽ|!��iy�<����aFL2��t?^�ogC�	�4�u:�D�.�[�͕���� H�y7@D�O�' ��@�Ә��ml}�8L�A���
���81"�#:�SSu��u�	�O����$�u��A������k���y��o7����y��o7����y��o7����~�_������~�_������~�]�`gC���t:�C���t:�```````gC���t:�@``````````````````gC���t:�C���t:�C���t:�C���t:�����~�_�כ���~�^o0�gRs�h(s����q��o�a10Xk�M�$��Pi��u:�I�*W)�?���k�'}?^�� eBi�O @��"�p��t�6��CM�;PhK���HH�u���BB!�P0��J��v:�(	q�H��n��4)t	8]O

����(L�)j����@�9�zCzC�ͳ-�Ņ�~HkEXWE5d���\DF�~#�$G�?,��^W^_/	j|��U��!�.�ɮԭLd�u �8D^·��&�u:�		���BD�/�f�'�̐��u:��B��R�;�T����4js����#���o� d՗K���t<��7@I���A��y�?]0a'��5��q��n7���y��o7����y��o7����y��o�����~�_������~�_������t:�C���t:�C��HHH�t:�C���t:�C���~�_������~�_������~�_������~�_����� �y���b��J0K�(K����H�y��o7��%�" �2�4�i#?���a��,TP8ۅ�^�O,�,�}�9���0��j�*
Ϸ������Bk%g_h9C$U3~�]�```g�080�E��dJ�@ꕮ�;v�65"�3���H�u=7F����ǥ���Xsi�"��"� �8	�������>G�f�L�O�>��8�>�)>'��b�% � ��A�K��E\�_��DTem$t��ۨ��H�]C}:�O���i�&�$$$$t:��#�I� �$8��` �A'��I��$�3#���M`o�4G0p�yB��(4��^nf�D���0w�A��~��]hi��w�K���������������������`���7����y��o7����y��o7����~�_������~�_������$~�_������~�_������y��o7����y��o7����  u<���FD���A��y� E�`@f"ϧ@��s�A䠀�`T �NJ�۷�����%r3t��"(�*"O�!�;��HR�&�FjYp����9���w����~���03����gCy����\쳵��T{�����>U<��`bJ���#S��",�A�P��EH�p������%������}�6?8/�)�n�#fh��0|>F#>.��Ha�dY�]�d�D����$İ̳��z�z~���N`�C���t:����H�{9:�7�����LA̒��2��:�B_�S���j��P��4=9���a%���7C�@!��u>�l�"���p�X���q��_������?�������?�������?�n788888888888888888888888888;���y��o7���H�y��o7����y��o7����q��n7���q��n7���u��n7�0��u7^O�����#���~���.�H 3�@H�Ҩ� �~���?��/#1{��^D8�Nwӌ�8]��"��Þ�ڌ�_��ׅKR����.s��΀ pw����~�I]O&��uEDA)��*у\�k�����7�!�C�!$�f4��.E_1=*��.�D8�5�  8�͏�	���`����@��)�#3!�Ad����Jb�Y�p3�8L̟9�	~R��H !��)�;ɋ���/���* o�`rGC���~��o1;�]%�� y��ĕ�N�v��P0�W��`�3��4��u���>٣��R�j"3��"	�*�?�Ĕ�7S�ĕ��CNC	��=������������������������?����������q��n7���q��n7���u>�F���������������������������������n7���q��n7���q����������]o����=�]a$^e��7�0��HHL�\XH@9�^�:)M)gR
�0��ɰ�9��:��O�W����� ^,���@��44>� �pA;J��@88;���~�D�O�&��6tV�@��}jd�TB�p���_�7�S̹��)|������Nb��wC�֒� }�p}����O���")>y2T<��G�EY<|0������RGO�p x��> �3�P�<|���(o5oj~�>�F��`�a���ӓ� ���C]b��C���y��`��@c����{��:��VI�Y�'갘s���mxVs���Q�R����Co�S�ݕ��~�/�>F�/�[�����{<�Q���@@@@@@@@@@@@@@@A����?�������?������   �q��n7���q�8�n7���q����������:�B@`ΠC'P �8s��M���GP={��=�?_  �# �y��$*��s��^^�, �Q �pBB&��K�]�h4\���%*\T�	@ 	�, �)450^Ae|�����]Fe/010 gS����pZ[�)�'�b��s�Gp��rs:\d��W'C���|���
(��`���'p~8�-��fY��D���,�}�|\O�ĢF?�
)����aq���FA�:�`H?�,(G�F�Y��u=¾IlWb�T��"�� H��f�}��$��#6Q ��0 0���8���[Q�e ��!�hV)V~���%+�-�0��A�4� ���U	)Gs9��@�g@�����iz/
J��5?�䇠�   !�� ���[��@        ��y������ ���" ������������ u:�N�����?�������?�������?�������?�������?���X9!#�0%� �y���	<�B\"�"A���;��, ".���b�1.CL�XzO&(�ӡQ��
u��>���:�\�m֣4R��c$�ך�[SY�u� �J�D9^X9j t�_��i.a0p@ �[���>]M����dc�%.�b8��.2�wK���~�rBDUn�=�TD�I�(horo�TT��f�e�|O��� ���'�S����~8����3!!��QfH�-�3 �m�f!�2(��"%	IƬ Jf/v���u�'�7I���&�X< UAVq�:D�COa���	IjiIeP}(��n�Ӆ@���4zt�\*�o��2��M���n��!�PH�-O �t��`@�8;͵@0X4L��4�5�"H�q�����Ā        ���������v�mx�!dM�� u���� G��������q��������?�b �   ��pa ��[�1��%q�Q@��S�Dۢ"�p���ĄBXC��Az�#Z�99J�*!�CyH9x!�!��s�0hE��^�z�))Wes������Ձ�.g��h5�H�=%u=�C_�2G;��t�	�4� ?��3 ��lV��Q��xh�1a7A��W8Ctݵ=��6���Ã L[
$B# ��f)(�>��>�p'���}G�}G�>'�.�Y@��}b�>�:>��&N2|O�Ap#�#�[pG����G��� s���K,�����L��J\��`��#4D�ӌE�,� y�������Y���n��$�=����t��`ʎ�5ew#�� �
^�	y<,��\�����1s� �8E�!��}+#����\n2���17ӡ�.�q�=��               ��2F�A�RK���q��������� ?����   #���                                        ����`������4W�#���fǳz���%�.�Pu	?C�ş�ቅ��E1�����\��� �J��c�E��d��n��	{ :_@��Pw��ӨI��y<�NttG���d�.LE��u�?�N0p�':����C�Irg�`�*�$��/}�8D�ۯ3�S��&��\�|�e]`����E�h������>���~��,��̂�dY#υ�e�8_�#r̜ �V�)�"7��YXAN&CZÓ87���$)C�Y��eAr�+υY�����s9�o�G���u����� �g�w�P��c�]����jYjy:�����1�$�Ϊ�&"�n�	=3���?ś��('
J�c���gls��E����nSu�H�h��u��`Ā��wX���.u��n�[���u��n�[���$~��^M'������    ?�n�[� ��?���[���u��n�[���u��n�       [���u��n�[���u��n�[���u��n��[��\��Ot��%J
��Du�=�/'0���Ue��]}��^j�"�\ot�I� �9��	2\����u���=���:\i/i��J�C��@��JH"^$ �y��QZ�B o�E8s�0A��}��\�N&��$Vt|c��⎿�`�7�;�@������t���Nc"or�aMF��6�Y	�#h��f͍�,�h�����
����!�k(��O�)���d̘�98�a��(��S�:��b�Η����+��� ���@���D��\d�$ t8���^�o�g:B�lxfβ �u��Ņ�F�%.v��K�K����}��8�^�M����#�0%��r${ 8����� �WC���).%	8�n�[���u��@n�R�;`�����	�       :�n�   @@X``c��    ����>ߡ'���!�Q'$wr�s��M� �y�����C�߫A�����%C2
��/T��b�1y?��	T�<���B/v��{���R�"���{��/�P��c��� �T.y2�_��K�� �y9�L���PP��n�«���R�VUD����4�	����D_O�o��c W�+��d��!��D|J|>|H��"��B(	�H�2T��S�||����8�L�>'.�[6�O����}c���> �4</�J|��|�/ѣ@'�؅K����1	|���ۮw��� f�(��·[��z $�	���O�˥�jq8�9�\�0dB���� ��|��6,�3�������,��#(�+=�]e���2q��cuY�H@�4�=.{��BB_���-�7�(c�$$$$$$$$00000000�� �� y�=�n�  �� �u��a!!!!!!!!!!!!!!!!��������!!!!!!!!!!!!!!!!!!!!!!!!!�!�� jā�s�B�!�-E�.7饝X8E��$�:�h{&N� �!� �
\�@\ŋ�P0���	��"�G�`�����}7������A�[��g��!��t�4����9<�`�C@�@8����"�|��NC�� =+�W;�u�� �S�̮� }�"<9���ܜ��� �������1>������,�&N2\�E p�|ҁ�x����(($p��*|���G�pY���0�#���ϳ�G�	#��l	=��������m0RW���CɕTH���y� :_/�ی1�R��u� ���O	,�i ��T��A���nY��M�J�zBoW|�7��56*��Q�]	�C^O�%WC���p������7��S�����$}���2G�ps�� �$ ��BBBBBBBBBBBBBBBBOL�^�A�Aߠ/��p ````````H``c��� t� ���BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB@^Ꭰ�Ȑ`0����� \�:ڛRDI`jϥ@0Ca ����b�"�H�^.MJ�kKt4y�r�p��l��Ǜ���d� ,$����{"�����N�A+��bJ�t�������S���x��~�  �F�B����`[Ow,���a0Eu��w��{�}�19RJ�\^�.�?RCpQd,*�db���?��!�Y�����!�ļh����n��ވ��0aaAAA5og^aG3H��*�HVݭcRA�s���3p�?��  ��O�w�ɤ���/VI=mg9#,�l�¹sZJu%��G>'�g��ɀ�f���1�b����R��.DnF�+/a�"�$G��A��An"@@G�������ps��,^�b� �����������������'���A�M�.�										u��d�� ��[���u��_��/���� ���?ˋ��C @@@@@@@@@@@@@@@@BBBBBBBB_����E�L�RLD`%�(l�F�aw��#��1�3�iY|!QE���G�ŀTR��=�K�1H��d BT�.����L܏�Y]/`��P30�gرW�����{%% $%}�����.��	K�AK��� ����L�:ի]�؎L��rxz�����;Qu#:ɑ�\�����,�(�Q�.	B����n�S�P�&(H����	�f��H|N��6���h�E�-�#�F�N���e\J�*�1��؊Q$n���a0��`��œ ����E�o�@s5� �[2����jrYi0#�og2�&�%s��� Ɗ' �D�y�(�Ņ�(=��L��֎ބh������.�zq�����P���rW��\��(c���u��?�]� %�1 GZ�5��0@�gSi�� �< ���J����I]a!/�`p���X���{�Å�B@^���w���,., �			TJ10T��KҐy=<���S(��R �U��@���Q��@���2�eeF,S���'8��3$�6b�g[���p�8_(�of�;��H&�1y67D�N���"`�.��;�X��$$�}>����'�嘦\Yj��vX�����������$�Qx��5�^ �E\	�H�z����/�|�5���p �d�%�;d�	����(��2p��y�,�>��p�#�|�(_�1�QpC�b|O�zDh:��0�p��a�.�b�ꡉp 0 ��A��{?A�L�����$Ot?�hb�OՖB��ʸ�;`��6x�x>ٰ����s�X":�x8|�R��X�HͩTi��dk/g	�*K�3������~�=�O����^�C}�=�`/qG��0T�PGP����.�����]o�sF���9�K�$881��u�ą���Ǡ�Q�{�����y��5<�_�!���p�s�$8$��%������������������������%����SɓTTJ���ȩ��XP�bTd���4biW.R�`{�:E�E�J�J�B� HJ^\�y���?��˓.\�S�E�R���h� �u��/�3����^�e���/���9��{>����ses�Y����we��rxZ��@���J�"�~���ҭ.1=p��p�������#���g�|�}R�W#��'��[���\�_��CŒ� �l��2fbPH��d̑�?����ܑ�bɏ��oaB+/��Ѣ�ǖ�R(�\�]��:�.�S���{��<ˌ��	N�*�������;C���|�4��M�M�Ě����f��,^�L�e����BR�" n����#!�$,\���y�,��� #�������Y��A�ʧ���a�`�r�0�#�Y��u:�B��_��׹ �q){�@ ��\�{��\`�%������h1��	/	 u��ő��`qrW����{���w����{���w����{���r����b�w����J��UJz�3CҢ���A�å��v$'>F��I ����zU,X�L�Rs���P��v�(b�gP���y����^��o����n�L\m�Ot:L����!��ΰ�P $w���Sv��jjң�db�%X�FX{d��y��ߡ�0%%�ʣ����O��̪�-����--J��J�nb���E���v�c7�֗���Ɨ���ƄDTtD%�T0Ix�#��muih�Ɋ��!����k�/� ��³*��K��zd\d�}��7@C�ʻ�}��1{�=�D\�@͈��7�(!)�ɜ��nb^�Hm. FF%% TZz$�$V?�=�@�/ ��2�+��� H�xey�������-���\���}>BOB����  !�uGR�hҺ�8a踀  � �%�J�y���d�O�����Oy�I�"A�e�/�RP�H�)(;��.^J�{���w����{���w���,,,�����S�^�0�S��d�%���ŝMH��G�S�p�8��dɽÕ§�=ӓ��:(U�ѤeC��b��.�biXbnf� Ց'S�Y���� )hs�*=��/��s7��!�$�% s+��Y1�@c���'����K-JM���a�D�4g�!*0�j�d`�Fי*ɁɂC[	�!�p_��Ŭݬ�	��֎�����~n�1�4p�!���0d8,ق	��P�bGًpqC�����1x8Cꦤ{��������]Ng��0Y��U1 .% / + ����O ŉ��Ϸ��u���	~���f����!�s���֐u��`$u���h$f�dΧ��"G����.4� �}9ތۯ��k�	���QQ .�>��ۢ�����q'��'���E�ܸh��`'�{��"�$���7J ��� �u�:�����/�'�	y���hD�P��$,,,,,,,,\\,Jbz�QO1Q]�%	���X�2��s�X���gn̃��,��OC&��OZT�Te�1c�����X�J�y� �?TN���_bʏ�w���c���`���@	���.�t��fA��GlR�/{�vX`��S%
��(����z�u# >�!-$����Q���3$p�Ϝ� GL�E��Ɋz�a���8!�3���[�p�'�8�8>PH��8O��8C��S4̇����qH^Blt�À�@`BTÝ,��5.������?�`D7@8��$�2u�CA� I@A�E*�oc�u������	�$��<hA�"�y (��A��&����
S'�
�17��km+9�l�ۙ�4H � }�_��A�#DTp�'ɻX�HKܸH0�J��%}'�+!4���rQd2Gp�����t���h`oaS��r�}�p��V_.8p�1�����$t?����g	y�+���%%./u�*(���ő�(�FJ ���P�IHNR&UI��.�. NO�&@)�XT�*�=^8��+��C���o�"�'P��`BT7��9��mD?���^��7[����H�n��0):0��1X�ŝ�:իH�=$�9�o�w[�P)x1zPbq����Y�E�'Ƞ�Y��Y��8*G���-�A>%����H�,�
"���> ����������n[�A��)�~O��*�O��ɣ��;��laH1
\�N5+�LL�@01Y]����f��P
.db\�p���O���Vghrs���	u��o`"@g3k��Y����,8-,�� ;�	�%�#�'J�Pi����4�$rr��ؒ�8_@a  �J�ꬭ�i((�`D��a"!�.�[��"�y��:�Z�eKΧCu<Łb��KP	�8ИI#t4�X)y�g'ڸ������~��I^�!��d�0����J�,,,,,,,,,,,,,,,,JJJJJJJJ�^,�%/
�,��L�j�D������bzzUǯ�A(�H��\ H��*`�R�bYi�a�)T�(���	=������?�j�� !��rG8�T�g�t�\!��}4���?\o��W[�\%�$�ŋpQKA�LcF;q�&�U<I�^�{�b\.��rW���P�0��CS�: ����6��QaAAD_h9mm<@IA<oWD7W7GGDV}��3�*��,5�� ��2�>��KD���I��4����!��+���s"4��W�^�7��2���d.d�b�H��u8�VP���O�ag� �5��ory�]N��I��j�R��������8��A�l���\� c	��T�dA�p``�p!�tW��W������NNy���8�A��D��BDPU���UK̞o�EGC��1� 7�����.,�.u��F�I�Q�^� @� 7�����H�% C�./=%��������������&ddD]=pQ�\@*��ϑ#������D�ӓ���.��x�X@�@����K& ^ zJ�$tҪx��U����}��KĀkAJ� Ė^e"G�7��4����fJYn.dU��1b8�,���S�s:��$�_�����J.zu8�W2)��y�m�Q(�\�@�"��J�R�˓j�����f_�d���͔/�ɚ��-�-�#2��˂~f��B��2�=ʼ�^ɫ�-R(S��!u�T7�����8��^�.rF ��i䮱��3�Ҫx�}�'��9ƚ��]/��;c�M��{���`��A����4dJ�
��0P�S�IE��"��.)��1IAaYJ�}��*���4CGKi��֪��O1C{��>��ϱSk�t����i|� L�_�.��Tb�b��#W���.�/~� ���hl2��H���Hh��4$��.�J\\�{����........%%%%%%%%%.�˕ł^`��#��-Z���:�LBS��̋�� *�������!K�*�P�d�DD�G�!ʄ�F&/�����Y��zz��d4>���F��] �Nc���H��K��ӥ-H��Q��\ ɥ�;,0���T�''�?�����J�\�MD�8����>L�|�"ߐ���@��͜�p6iy���R�ߖl�"ى(,�����EY���c����Y�m�"7d��ƒYY�^͍ ji�-��E'�=�G���ZD��_a ^��@�N`�q17����Ь�3r)q�@�bBaL�O!`��Њ#@k���t �6>[��v�`EE��0����f��?$���
d�Rz� =}���	���?[��B���J�J��$��gs�'��/��,��"8����Q���&&"�/�g��X�81�&�%FOT*�	u���>�BA�G��D�uAgZqЗ躉(c������������������\bJ� 2/	�!�3ܹD�9J�%�	���� =���Y� ��r��Ng�2�`��yx�̑D@�)���R�T$����	@��.F"�g�D���IA`@�Ǜ����� �}��JAM���Ms���p�d�h���,�0T�ң�� ��'1v����թ��2sC�h>ܟa��fAl��#���&8�	�pL��ߖL�N	~>|H�#��|�pC�>�8'��\�_�
H�z�2G����+�����\'F&> M�Q�2�2b/a%����.�	p��.*�	�:(
�a���7��5��.�����=�9<��0����v�WHI����{�q7K� ���~$Bt��&y>џ·��8\E|IpqqФ�ѡ 01��EV��qqO��`�rG�"�А��;K�L�%�$�X89�J^b��\ �.u�=��6�A��=	u�:@�^o���� \0E��//
�$F.................../%  N{�GNO ���<(�(i�ck���s�R��A�V����A�%�硢⎞��TN*��qp
sj��穑���p @�.�#�Tf ��bS�	���0K��81\��L\�g_jH8�,!�d��@���N3����Yj`��L�.�5�JPV8�ɹ��.r�mhG���~\J�膬�! �x�������m�eA�%A}]��	���r���s����?ߩζ�"���$.�.Q L���'�0s�=���ju�?��Ā@��� @�%`����c���|��@�.b�W�`�@x�����n�62���
Ws=���&:�z��<��������!΂\d"�� �s�#��3�=�".�c�BA��A�Y_BD��5&Uw@�H�k�(��t ��J^�$}��(�'���D�-N�P���y�8] #E.�C��J�s�����VD�K��׻����������������q(�qs��&^^A*��y���d�E0*9e˘�JU֜d���d�y��m\)(�rg�s��K��	Rj���B	�I[�O'��ܹ=��M1 {�* ������7�Ѡ�A�	A�@�� 1D98b�`w@:��Yh�q���Yjb
)�$� )��K.�RlK):���E��}: �"ᎂG�����p���/@Bbb!�BBo'�Dh 48	�}$�ٽ ��]a`i�]Y���"�Yp��`�b�r�b	@�e��{����>_��g�;���IY}��$j$T 3jy�����fW�0�(c�ֆ�Yy	��%`V4	gg$_6u'�=�B�[��e�g�3���\ҲJ�.QTt��",�� SC��Hh4�.z��}	��/a7�3���j6jh|�/�^��HeK�LC�Nr��@[�@i̒&���{��F���^�� �����.��_�e�����Xa��������yyyyyyyy�(�r+����2 .C �  ,��Rޥ��w bTYDY=)�+����7[�qI��T����˅TFv@����bz^�C\b.� u<��IA�n�ۡ���}4�A����7���AQ����R(�� ��\"Р� OKv0���-LuQ9<)dde.ɰLtQ �J� ����%��v�cTsv�?�@��[!�f��ct����ܿ/�p�۔r�-�nZ��#Q�uvB����q5ihA��:D�-Od����&��:��E9��#����G�`0�]� H�TO}�:ӟ(J���	$�����  � �^�o�3�0 Ө�TY�i��)t��1t  ��� J��Ǣ(�coN�(c�X!�4��l��t��:ϗ��\�%��},����_ O����#b��u��
?H.O{�?�P̌^�Nq�ׄ ���sF��23�P����)�s�5��{6�<>�������$�b�秧��������������'���e�ε�{��9����2�'*�J�Ɉ ������t�Q�Z�:bG��=3��H����Z�4&���$~���A��#'
	)1}�99�@�'�**�Y����L�n�0��a#M�3"��p���,�2S$�2D�X�*:A=P��PAd� �
HHq!*�8���B��C�EH��2�/�Ģ~?���|AN4�Ȇ�"�����Q>�� ��
HIK9��͕��i�&��c\1�b�K��f �C����~�6��ΰta`�g�0�@��{�
FV~Q�Ϥ��`Q pǁ���s��N\O !��1���1���9�^X�����ϣ79�(hH��0�HM%�@���@�	yy��}����!>[
D�ncG0���,�jp�"���4,#���ĄF�Ġ'iX	_����/���4̹D��4f^,\�%JbM��# ����X�>�fo 	�@C�L�BP���������LLLLLLLK���OLU˞`$���œ�P�ov*!]ݻ,�ę2Q�$��'���C1`Z�)s��;n�T%c�(�I� �=��GH:`p�0'3�)p�Ȣ/r����:��������$n��^�0��J@9�z�M*�KFFvXae���{��FTJ����*�b���N#�"��>��69�_�p6a(d��zP�m����l�p���	�̳�̾/�������&a#τ�f����~n�O�H��i�rފ�R�Ĳ�k�FCR��%XX%Oy:����@$��Q�ӄI<DY���ln�� J^�U�f.$�}�+�����c���E�J�O)dz���&d0���Hz��&"�P}�L���HBs�)`��7���.Doy����=�Sŋ�Ɯ�&b�$�O�������֐��d�s:���OI_�4eG��`J��y{�HUC"��@��G0���L ʹ%��}:]	��_`�%�j��(hhf'�ĥ��f%ħ�&%秥�j�%ĥ��(e�,
���	(剋���Z(t���I��4�!K�=*(	Ɋ�6	`a!GB�
u��\�㗅�s�7S����OCy�QR�t�� ���J�1��^����d��D� K�O�wjQ��1(�ݖv:�+��Ā
�CJA1x�ܹD�X��A���[ZCx
��(8}��PH�0��&b�3GĎ3LP���~d�s�UTCDD�����3Bʳ�ä5����Ù��F L�r�낗*T	y9��m�t�Χ�J0b��Y�"��.�u:��N&Wȹs���e)3y�� V��(+��/s,7T`�b�o !�pG����RR����Ǐ�QRΖ���ɢ	�C܀rr�c'0���#�AE����m|������=7�:�n�O�FU�����(�*��L�4���d�J�{���������F���b�.�<��%�%��O�6ѦǇH���5����*!��������0'�#(��!���!���*(�����XD)ө��c�Q��ĂF/`�ZQO��ʂ��.Z�0��Q�W)/L*�4�X��w�D	A$%��}�].���K��%��cD@*ך �+'���	CBb��^��	Ө�cK��gc�b�++���P�A9=Q�&�{�\�xg|����4�+���VW���\F	��#St&sDts�ĔtVv�6Vuw��̾��ξ���~0~�$�8�W�̄��K1,r����8��^M�qS����t�����=�o�%vvBBá�%��)4s/ 	��BKԉ!	�
XlXr9<Xm_gj1s6�����2!��}�'8ڀ����7�0�zs��ڼ�3s�* 4�\�"n��T`� Ƣ�����b H�7B_ey�����pƧ1�`��� �� )=ڛ�pc �����  b �~����I��2�

���H\��bdd������b\J^�����d������ddd����]D��=��J2a�e�%b�B��v�\�q���i@��	�1 �C�z�jZ� �\$A�$ z�t�ˉ�������]bb��p p�d��[U�	�?*�珧�H8K��L�X��H����,�wn�;k���. .Rz\�b�p�����\̮��ssDw6}�'��|C��#υ�2@��(H�H�8/���8EY���l���,�zP�ۓDW!x�e$��o6Gg|[і��:��]l/�q�K.{�%*�d=�z��P���^d�B���c�s��
q(66�{���$`u�����?VU�˜�	��ďH*��ș�0]=��&����U�`c�"�H
əp�J2�'Hh�u]|YT	�H�Y6Y@$Ey��TO.VYP��y2��BBB�����*��ʄ� �ǡ�l�n�@G��r�����)(`� c��P��u��PPVy ��*!�������////1CCCF1��TE����'�00*'^!R�F\��e+dœF1\�:�~�L��,��QQ�K.TQu=���J�h�'�%�$`f  �
L��~�����`@�
+L�j����J�2n�9=�Ch�e 2�ݱZ��2�Gv쳱ֱJ�q�BU�rS!b�Xhs�4	侄�RQ?!"����W��d7!�B�Y��f$Y�E�fH�O�Af$p�J�qd?,�6ܷɐl6��X5��F���U�L&���4W&�@�5��0b�e�TF&���L�]��.$~�ߤ��%!�%�p�g���@s�/����E�� �C�B[ ł$D��@�.���EV� ���H���8@�I�&�U1C��$�r�bbL��+�إ���L�}�"e���B/w�r�糙Ƭ �\��H0_xu(�%~������І�Qy C*��Ԟ�E�|�9D� �7��Q����0 #�� �EQ���QQ�T1qc�`�	����?�αc$�d��IɏKʥ1	%RT���Ȩ�+T�#Ա�NMOF
\�QZ.���Ԩf*$�&%1{���(�͙P_EǠg�e��{*u	���1.`OQ ��r$t	�����TA�b�1b�]�1JL��ݻ,�u�B�
�L�3݀��\�0EDŁH:��M�pC��D�"ٶh�8����b>�/�G�	�(,��$T�2b>�,�����"*|��PJds��[�F#>/��ܲ��B����nMh��	�r�jWFH'1Z� ^� :��O���4Xɡ�4H�{�Y]j�COMҒ���I{�	� �@y=̜-���U��u<��, �>�D[�b����"�T�\�$$^b�LY��F)u��x��1H� ��iU!�E�R$��QQV2 h.#�M����I�K.������g���� �#?�fz��]P X�Q8�&�	2FT=}����/��V)�OO_�qb�%���M��n�����������(����'��#(�����X�4�$��G
u12�E;�1'#8��:�^��XQFJt��lC��FBJ���`�A|&��\�^�N����:�R "��ˈ)�A��f�Irq���u��\�wn�;k5DaKW=Ɨ?�b� /����SQ�b|���� �n�B*�,��g PR�:>�#��>r*pH��d�Y#�4�/��~?��H�P}�f��G��f�wS'&UV� ''XU���2
T*�y�8c�Y�,�h^�1��"f/w�A�W�ȓ �P I#��$�z��$t��:��^Oײ9�5�|@Xi����:�B~�)z//O*(���f�40�
���c�(�hQ�0G����d�4\��}�x}��ZA�L�C	[K���H�/G�w�HX��Xş�` `'����r�=JA�E|�72T.{�����@߯r纫H��P{����dd��(*z踸���ps�$@0���E8�S��0�'����b �da�eWVݩ�,X�����F/��s&'���N�!O`�  ����s�U��{���Y�zM9)��a6GLQ�]a��T�,0����c��X!�����Q\��V#�vY��X��%v(%ԙ��2L�L�~��^OAa07HӅ��xx|�Ş�כ���}>�O��A��=�Co� w[���=y�?�O�����n�	�,6�5�57@�_B�K���Jz�M*�� pg%���
s�DE��q�?\�G��4��	&^�u���� R���V��/��"��K���{��۠�/7���Rd�$Z��ӫ��=s�Sц�����L_�����3���i� !��@���E�H#�� ,^^�}�,�:�\#Nw�����69ğ�ҭ&�j�� ��W�Ӭ19�� j|�)o/�z,�q�˃�D�&�����������}<��I����0U��= 2O~�
��������Jz�Tg���^��z3d�0㭮Q�J�l��R�,�8�閝`*8qqV�X���?��B�=��ɶ�
^�~��������* �,d�n���m�6hm�X�9��h{�� FCy���:d0aԤ�v쳱ֱzd���y�)ဉ��b�0�q6v�3uΠ��|�6���B-��b����S���ē�vƅTS��֮�n�`qq<9�����!���y��y}��$�q��B�ݱR���t�R�N���?JCJN^a�3Ӆ��FCYs0
{�:Q�N���o%�tG�ä���0��#'���qxDk1
b�YQAr.L:�wYzd���n��:*�/��47���)rf'��@@���s2������ī(�����s�Y��hru��[LJz,�����u��̕�����@K�X�\�$�}����l�D��!g�� �ƨ 4H,J^(�  Jbbd��@Rr��2�e����*d�U���/ZU�����)x WkS&[�R	qE��'�L���2r��K��:�)�AW8DK&=x �\�T�1袡�@��bW��33�� @5��)?�8�W�����0��!�
�=��K
Z�&�,Xabíb�A)V �K0�=s+�T~�����
��@}��C�C�pAF�L��'�p*E�dx���Y�Y��p��[2P���o�,&�	ܯ*����+9!+���!?@�ۯ�q���ݦ� 19=qd����D2D�Qg؈3�Y���:�B�L�#j�h�� � �at7A��EP1�,@8!�7p���\��7ؚ��(s�@	����y:ʥt�Q`��!b��(�-�� O`�E���Χ�"oqbWSS�=��}'�<�(�� n��Z
A�	s���EŐ�ņ%IrT2p�!�� ���
�� h�8*y*{��P��逩�3��\� �i�'SkCu��~�]e�J)�''O2L�P��S� �8�@`*$�J:b��:biS1rV.֣�̈
`
�14�L���:�d^���S��b�T8RpH�gd TQ��������Ҫ��t6�<�_��m��T6�x89���ܖM���J�����b��b�)TɎ�*�о�u?�d��0WB�
��z����"߄�n
%��b0(�|/��8�,ӂ}�������G��1"�&pL$YAp[��p\B8��
ex)q�XO����x�/v1s�e���J��^du3pI1w���β ����d�0gӤA��&z����-��)OL��"��'[��D��&n�E����a��'9�P����b�$��F]{�8�O_��V����}>��� ��L� �C*����r��	D��α���%�7�#����hҰ���.:mPX� �?}�9�ޜ�B���H�/p�ѫ���	 	n���Ð�Sŝ$�.س�!X�4&�n���Ƃ�a����H

+1H�I��&(+1�ܪ�A����I�. �Ls��EI]aæ �^� 
&����U+�̒�p��BG�qx��-h�r����GFu���ĝC@���b���IeCǑg�������2ZH�}��/�Z�*�Ɋ�۷c�\�ĽDQ�*\m��p���d�Յ�2�CCz���&f,����٣��J<�l��#�|��R�pH�~�>wp3�"�|���$p��e���p_�ل�����pܑa�"��ŴP��;�pY��.0��%��
`���vA==*�g�" �o %g;�s�D�E�.�y8�J���� ҁ��x�0K�M� "���s�"%�(d�S#���m_	:�j ��3ع(�@��� i��.�B@A�λJ�s�� b�z��E� �Chq�N}>���u�T���#���� �.��;C���r~��bG+*eeW�t�C$g�ps�4 ����y���0�7˘ !��q� b/  ��'q�pQD�OO*U(U��3B����ݮ:���<��R�2���d��L��AYzq5!S.wZ��P9hQ&b �	 X�U%�t�C���n6��	���d��!�����˩k ����\L+�8���I�L�)�u�S)*�z\d���1��~��`��!�>ۄ��٩|/����,�d���'��	>N�N�H����pa8�8$[�fȶL̂��/��
0kod�żݺ��`�R��А��\�āi��bU=���"J &��Z (!E�z&�f��q�8��6R$�${�TbN@�� �X2	40u?�?[����u⑋����h�^���4����Ġ*�p; è�FH����x.Q`{�<<�
B�����+�'��0�ˡD��R�"����[k�3�H�U��p��9?�	Q�fD���tat`����ڰ�n��u���E��ׁ�4�P�bb/a �s%��0'�JTQT�3$46$��PԪ'%2OJ�����\�D�qb���F2u����v��)��NT=t ����*(�&u+ͬ\�QD�$\S�@%99HW�1����A�j�+�`O�<\X$1� ��])��:)�)3��8�X�R)�P��J��"���\/g3ӝ�x4���4R��n�ܚL�.��V�5Ȑ#���}	:�����`BP bG�`8�����}�4�<7_���)
f��e��8)�v�v'S.J�DX���+�Og�0r�됱���@0J����r�&�l���K��J^�FB����X��._$9#9�^�+].7�u� �R�Q\ �h)`��W��0�P�27Zrv:f+���1�4� ��M<8���BHhPWXzDB<u��&,�1d����T�7[I�':��.�7�ʠcP�ɥ��t��A˞积瘑#�@�f�}9���n�!g�1p���8�=99EQQE�QIE')`OT11Q:9)�˂�J�v���d 	S'���� .\X�RlW*	��'':u�f'I�R�0�s��\��%=&L��8M�$db ��*aOp�B��3����rt:�UD���J�� �O	/�
����tTH&۷c�\��QVg�c�!���	NLz�3}���BjA D�a�#COדkiI���Ύ��y52��!5�0��/�������7����Ү�s5=�ڞ䎢�ñ:q2�	��Zb�``?�(��_@�)U���U�w��� ��� t�	��,�`��7��J�/1%N^|_O7�9+�\D���TO=.$rA)u���F:�]@n���E=Ӆ�ł�\' ˖�3�xU@�Z�Ԩ�d�Qu�\1s�I�����xGj<UPn���ZĴa�EF3�!7�0��N�
\�b� �1gи���&$�`/	Ty<���[��&�YPp������?D��A:t�r�zq �$	���
 �d)JW��22y�5ɝ�c��c&�X2ҬN��J$=)�	�&,1��&��iN${ =�E1.NOhy���Z�\�1��t���ܕ��рa����ٙ���Zx����%J�\�b��b��$�C��*&O6wHc�̔\i��@I��50�����~Z�O���"�#2
Ha(!�|��~��Y��Y1���fi�d���!�Cȥ���]���l���s����*�J�/�t��d�ŋ��*)&��A9��t���� D\����8C;XC���H�Uy�~��>̏A�BN��K�M��t!��<�^�n2hb*�OАc������}
vLHȐ��#���7)v\�r$`:�2$}����
&�bd0���c�%@���b�'S�Qd�H1��.(�8�k'���B���A(�.p����A�ع��~�>���s�@0�w�A��������pL�-��g�.0G�p	(�H�P�T�0D�9E�$�\Us�S��LP�)T���\�T�U��ST��&%F;Q.TF.CR;�wc�\ŊT���0i�݂ ��Tx?ĞΧ�P�T_�D˃J� Ǜ�h84م�yaD@��� 1J�%�)�ia֎0`�X��X�J@(�eJ���_B )\Δ2���6�F8�!�,�l�Ͳ��ۆL|H���($p�Y3�_4"�ĢFpY'�G�׀��j���e`�>��I0s��>VDϭ�mu�W��������$Ny��Q{�$47}:��F`�
���0$�. � /u��!���_$E���i�G���_�J�D�Q�_e��*	U�V�;R��X��)QAϧ0��L�ђ�*��&d���s��%��u��W����=E9�O�[F=�u���`=%*�p��m**.�K��H�$1$_WHV=r2p��D���B@����'���
TN1
(�9<�1�i��C�P��U��s��:���1T��%&L�f'_�!a�V����T�De.�-�
�>��/LR�r�n��7�ap ��'�����O_`���� P6�X��A�T��}P� U)��"�]�L��b�c��c��؝L.x��{>�Q��fm��6�?��E��jPY���2�Qω8'ɒY��=d���,�A>vHl�q�ϲ>}��pC�*���hHcs����f�<3|�?��v1j�ɣrU+�
F����u�R �J�x8�4"$�>@��bw��s���Cy���F�����{�`�+͋��Dd Nn��<&q,�b0���#*@�P��%u֙��^� �\��r���C�2U�Ғ"�2%Fn�&
��C�.zO�Tt�����7S���/t�	�]-�c˄�u�w��"�u�,A�D�+���.QC=�����כ��QJ�.��C��UH�T��t�C�S-Jt�7rɓ;1r嫒���kTX	�����J�*r���s�����h�WR��R��?D�@�d����Rb ,���x}�92��(%%ɀ[
\%ˉaS�.b�ե��*�r�#;i�*J�T%TF=u�!��=!!(*�L��l�8[�0zP�����"����Y!BG��B�O��ωAf�l�β���
fۇ>�:p�|���&~�"�:|,,%Q2�w���JK@(�s�M��N
�2��V�`&��(�̒��N,�|��6   �����c�	)) ��)� �:u��NOO}�M"���o�,K�����I_O����g���{Z�(R�&��"�5bb�tR�Х���S��(dk�d�S�.2}*��4��>�	Sҋ�'���*?��E��2�{������e��!����� �t8B/��
HH�s�iY� \,)�1�,�	C��&EDQ�2�A w�sR�{��@��5�"D
��-��*S1\t��!���E�%ciɫT��Dg[����ΝJ�\�}�ұb�8�$��TGh~���1�r��"f�t2k톁$�NUB�2T�����,��ԧF0���G*rP�aa����b��r�|O�B" -�f�d�3���YA#̑�|Y31(_S6���b}�N!�p!�� �6�� �����+�9�Td�1\X���Ay'����Z:�H��W&bXs�R����8\"O��*�/�`�C��3�}����	~���>��ZAD$���5U��upWX��9�IL�I�]J�ā!�哕$Ψ�'.F-v�����dӝ� @���\.Xź$�F\@���46d=ˏC���S�E'>�*T��bL��$t �X�ė�@-BO ק˘��u:^��η�E�z� J�n�OB��v$�HL1Q=D(���% �(��3�2gI��`��'N1
M+���0�8��d�E%FbA9)T⤮�䫉���b���b�ِ��c�fE�A�!�kH''���v�u���� ��� m꤁�(O��葕%�hLi�(P	)�j]�N\�䩗),0`��ֱ��'_�.��H0�p�H9��t���D� �ȓ���8���b^z�UH��ybø�O�` #��H�>��BA�Kc�L�M�"��Fs>����rҨheV�\X�c�S˓�D[�a(d�R�^Dщ^�[��h��R�}?D����� �!��<�K��\ �� �J����%{#�?\��Ho�'ڳa*rf4�)C�N��*R�e��b�o�u/�d�B�
bd �|�+������j���kO_��1b��2���M��� �t��-כ�h5�f&,�z�~��_op���%��	�b@���t��	B�&���1 C��5���*�wd�&,�k�Lb:��X���.Q=`*k���XDɥb���rR�Nλ�t`#!HaE�FL
*'I���� ]n��0u��1�V�G� j�ˀ���:\a�7��!p3��*k�R�,�����,X��X�Z��x ��҆f��p����I].7;K�%a�a�\�@� L����|�F���g�����f�B�Ie��ք��@�YĈ6g$1&A1d�F%���n��Q�*lG:ddtv)�qQI�I��37�QP����� �H����P��:�@�Η�ps���	NN	�b�e�P%�b$�=�+<�����L��B��L�~���VZ��Њ� �s��i�.
��ș5�����
Os:�β��!e���2��%=����1ذ�s��P��rs�e��s,�	��5+�*=��_bF��`v�&� �`��``�@7�7�� H�t8���1�'��pq����M����ɡ��,���y3��[�R�Q����p�d�N`,ą*��q@��/�"P2C�D�&)s��Aw��P�
	H3���4�~�ĉ �]d���i#�9)�9s�j�4�Ŋ�,��vX�gc�\��91��%y��_Η0 �����9����%�x���	����$cSd�&�u�Du�C0¤˅�d��� �J��JKCKK9�i*2�g�ŞoeWS��v�YiTੇZŊ��H'(��e�/u@�� ����$B���ʮ� ����jH<t����_Ϸ�1(r�����	hn��\�C*��NN/  ����u�t�(�:�N��J���Q2`T%/!:B�<p�JQ�U��	^�7��X@�1ԱA�� ��ߥǯ!��UG�	��a���.^A|��]�蓙��~�:�o��1#���&�}!�:�B�D�`����99K�#$cЩ���H\u2�*��wybы]ӂ@\`	Q�d�1= �2d���*�+�LS��j���I�@Or��ѕ�� /��� P�;r��p����!G@��������v����ʋJ��rŇv�gkX�L1i �A��/��"ĭ�;���}
	Gq��К�^���	-.wP��u�e����3Py8_nN@�Φ�sv���`5 &��S�a���[t8]Q1q[j�2���5ԩ��QU�V�,�J��B�=Á�̔XSӉ�ī��D���K�+OO�����
��UeTR.b���t����/�S�R�(ɓ���6����֪**V�q�خR�)Х�����IpKCk�Z��;=ub\zd �UQ8Rz=K����rU� ���t@H$$5�\��],�.\J^�DX9y
	u��F�b���7�z���`N=`FN	/F$NR�H�u��R�Z�=�b��B,�u��*�u=Ej`�I�\Y)�ɉ�Y�bî�=T%1��P�i�1 �İ�xQΥ�M.2Qq�����Χ���j��X%$M��D�E��R��r9	q�*�?�T��=�HQ�����:8�حb�۲ŝ�b����F&KF����II艟%���qHi4UXA^XmlUxm}����^�F�7�C������ڐ��_zXW"2H	�Cm�[��\^���s<���.3Ыv5,	�؏b�p鉅Ct�^eL�E#���:^\�5}	2�((�>�/3 ��	���BW��p� �0���W���J��)P��@�!+���.u�ZLbe'Sv@H1���a�ʗ������)V�C=NFZ�� �u�'�J���E���/[�1|����p����w��0r1�2�2�����Y�H�h4ly���b��ΰa`�L����0������L@����`��A�@E
T���K�EZ�r�E��ܩz���S&9ӫl&WkI��-v����z^�F8C\a��.��A  @��p'	�J���H���%aEe�4�B�TI�0; WQFZ;�n�Z�3�n�jի���t�v�}�	��HneG�
S�|�QA@HnLי�/�W���Lͩ��y: ��H�! ��XMd���jԞ���ͺ
�8��N}�oWok_it���F��ׇ�����q��m�aE�?E���C�ӕo��CK�X��^`�
Π�Pk��"�&b �% y����o��p����Ȑ0�,���Q�I�H�R�+A�1�q�d�k��Η%Z���ԧ��2y��J�\0�re�Ó2��Ë��:���O�'C�:L�c�EC!�!7�9��Q����*)Q��F2$p�0F%}:���f�AW��`qps�D�P9�&z�u�'%F��- ���/&�)A`��k����%&���tRqU�V�F;qݻ�/{���b��gkEY9�S�%��FO
:{�P(��A���}��߯�g���q�� 
ʭO�� ��D�mAk/�QJ�ӍQ�H"&�cK\�t�J#�vX��خv��㎵h������ ?�!d�_�L�������n_�S�~8���\�-+�Ff`B/J)&����,�3[c**���k������6�j�oq+�*�9ޚ^mѡ��0�c�\Y�nt��Ԯ�ZV�=�b�3#ҧ�0��d2�)J���3��:� �/�Pk��Ju�Dɀ8M�f�z�T%�\�u)�`DaD�5Ef�  G���t_�r�& �+�$�5F+]�����\^.�q���v��y��1ؿ�n΅JJL��4bdR*�`2u������ �)6g=��n��
E:ƞ���D�� �y�R����M�H"�}Q		4�\a�b��L���'���:��))ԣب�?K��&�A�1JS
:0bT�W--��T=QT{ر�:���bq��LI������= �����/���$Y%�b��f�t:��@�ba�קS٩��/.Nq��@܃_�!�7�d��T�bU8��Y��]�v�q�ZX����)J�L\�ƢX 0+�X���~�:	�7���mlt�����g���. ��@ 9���T�4f�%
�C%F`F&(X\� ����$�	=O��0'�\�۱�Fb�9��*pJ1���d���������$�p��������aX� �
�u��''�
Qu�RT*�(K�I�Ń�O� �� �®T����+�d�����N�.JX������vĲ��f/2	��,��.C/%~���/��@w���,�bT�$����p��+�% !��V|�ł� 8]O���0���8"� '�����$Dt��qd7��   z\���RUIgn�qT�7�z���b�j�k�S�1CO:>1��TQ�`vU,��ܔ��t��ɱ�''��=`
A(S%�J�$	%C{�αC$)gPPeq�� 9�a.�c!t�ȸH��j}<��	�B��NZYk��,3Y�b�ݻq�v�h���Z�Q(��_եwn��iG�AD�/�`	y��<Ã�  ����h��%�"�YeEg?�$C��!������ѕ��Ys����-v)�ܵ�ڕ�TV�^� J&�1��9��1O�8P��S�� �n�����=$=R����	12,��c�9��/	NC:@hh�����rQ"&����;�*7wLz)l`�L)qe9*zT�o�@�4��LOLDP��3�g�yt4��b�(d��&��qd0�@B�@��.07�R �6�u=����A�'��`O7X��)1p��"�ǘ�  `3�P���%N:L��æ\�1RdʐJ��e�Hĳ���J�w�\�c'TIK@�gi窇H;�R��4ɇ�c=q����G=�D\����.����˞�"-ӒG�K����q��AbN��I���x���t	�%2���ib�]��,X��n��gn�rє���I_�ZU_����7Jʨ���% ~���D���a�dD��b��'2"*�Y���U��4�~_V�sG4
k6q:A��` Ґ�˨���R����r�����D�H���d�|�(��]t�MO��8������=2C	O1t��� ^�X8��z @0A��u{������ġW:����k��S1JyqV%�1:�z,@t�L Σ�㥊���1.0��(�?�o�!�d��N�Ë	��Q*�β�.����`�庠���}���7@���X�00�Qc$���p�%��Q=Q8�u'V�(�f+��L�2TÎ������:X�����n�L�T�L�3*a��K\=hQR�  @r���M�BQ����L�V�9��/���4�'  �5;���%��Q�L] �	�Lt����n0`�ŋ;v��bŋ,X�b
,E1�fD���MMM��/N����C�5��4��$�r_BA?�(OO�B!�Pj��m��zp���ZUO-ce�����5igd$���ڕ����Z��˫Xئv���Hs���&z���H�
^z)D<~�" �. \�r��J^�T��T}��~����#����Ft�	�\zT�-1z0�jab��k��,u�(��K����ewY��S'Puj�r��ިz�$y	*�ы�ֻQ{�Ft��M����#��rE9IEs�8���,�$���W)
d\�T ������..��*U���Z[L�U*T�Lt�T�]�� �j���wc9gc1��reɔ�L�r��5+�;� tv5@� 0@�e�A��J�*R�V�<�o0����p�� �����OCb\J "�y����-`ZYqR�X�Z�wc1�,X��n��RS:��N�|��X�R@�D��ۨ�� א��H	A]���rΪ��y����]*�Ow�����e�����QkH0q[�i�d��	A8��H��@�I�4UH�����&Mj�XX�=�9�zŋ�}%$\i�AH{:�E��hhi� ���b�@��������]Nǻ��1di<���^z��.ip�

�J�HH�* �(�1gc�v[vu�P��9J�,E̶ A1f  ���aeA3թ�$��ηC��� A8(I*�`�d� ��e�WXV+��2JĨRQ6��~i��d��,.��{'��%Z�r��������ŔE)q;�GLA98Q��KF1L=�V%���}i�JV�RZ1�(喩
.,�SҤ�.ZX����d� ���(
rT���0�B���3 ��C�G��/�r@v/g���h#�$I���CJ^Y� �qرZ���0�gn��R��Ju�,&�Au��������W�7%����a��E��fC��hf�Fj��i#Fg',�-��'@��E�|i�0ad+��$YB|����p�"<��?(M�#AE�J�!�O�0*(�y��'� �I� RN��:
VF�.1;Ì��z4���^(����z^&d�C�u����)T=<s�:W�
��*��s�5N�X�ѣ�`\0zҪGk��kC ���HkH>ؗ?�����T@C��, !�����/y��!� ����ZT�2�a��M� J�J�t=��K��KԓQ\���.\�)q�cC%�*\�;.咰V�*t��p�X�R�2dɖ��*CL-���R�2%bu���s��K�ƴa����E�(�Sb��1s�*�]"�������Ur}��A��:�bB	���0�S䫔�b;#�:�r��íZ;��2�ӥ����P�F�^���iż>������ȏ gʻ{ ��&���
Ɖe ����3���F��x�t���JB�Mf���芢�r�8��Z�����
\ -�I5��W
=
Y��Ja��Ү�	cLT��DL���ޠhjt��Y[D_N�C�5 �`�A����Z����4�"��C�ΖL(��"�2R�t\Ȫ��d�ۜ�u0H�jqk�H�ūJ�1,8�"�=����O�@�gS��<��� J���1:���y:�@orG�re����X� L��r��9QɁD�STeBPj�$�MZ���UIT��I֥�/O*us�ũ�)R�q��1ֱ\�2eŇt�%0�U��2r��@��K��"����ʥ)+J�R1Jb�f ��e�Mp� JW���݈�k��!��F/T*�s7@����Q �2���خb�3��,�v,X�Z�j�,V�b���XD��H H�h��{��O�`������ ~����E+/�P��uU�6Z��u�mT����x��g|�������0�2��3�Q���f"�LXӕ#�b�D�Qɘ�R��Mh �V'V����E��Ucg�����.n��/���`ﰀp��� �}� ��ZT�\�Xĸ@1�����b	_AH#.`%S=3mT-\,)�S�F*��W2/NNQQFmjn���b)P�1Q=<+����ʃkS���2���>��d�l_b����"���� '���#t`QJT_�/� ��L�)U�KH*)J�q�q��gkSS#
 �rŇZ��a��JQֱ\�r�1��R��(��y�(f!�#�T*���R��`:�12թ�1&�ы�I K0#M A=�^,�dL�9��C~��C��Ӆ��_n�X`���Uíw�=Ie�S-s��u�0�grŶ$ɖ
�**Ar䣽Ɓ���(��J�{�06�:�M���ϴwx������%�8�^���pՓ0g9�"#2F44m<2+
�H�W{8��՟�� =O�9D)ҩ�X�Zd�����i�����@��8M���%���u?��	D���u��`17�pb1��p����ĕ<���B��J(�j{���AD4DV�Du�S�T�3�֮,�m�4ʆn�'��9x���Ą�r2�כ�k��$)�z�@�� �~�>�%ʄ�W^�B"@�s"Eį�;a#������u�N=&uJV$�.:IRɅ�ǩV�)J�b�i�;֩J�3�ū�G��V�X��d��\Ĳ�n˘�G�
�t���B�v0�r2��r�ةZAh��.�J���*"�iU�3�˅ :��D����-N� �0� 83�A@D��8%��U2f%��2J0s�V�L�s+X���b��h�a�,}�0`s��P�p8 q�p;���K��f�|�:M���� 
N�J�;;t@1�.b�d�|��,,�W����:��W܂_���T5I@�z{�R�����h�7ԴŖ��/= Cp��=t����� u� ����49���J��IWlT�RU8��x�� b12�C+�N�R�rpQ��F1TZ�P��q�1a4e���uka#Bn��""! �OqpGY�pb�9���L�X<8����=N2OJ��< %<�d�D��ӌ��vZ�h�gHZ��$��
S.,�J�%�*T�`��-�:�,V�쳲۱�Œ�b�u��R��k�X��tʂ��h�H\0{ .0'�T��&�1{�����Ty�:�QM���A �7K�XR��T�]��af*�F�*щ�&L�s)��*@*rs�˅
c��c$����C `J� �^.�t8��_n��!*ps��AԬ`�|�	�����n�$g���	�H�~��[U�&m*/'�����9"�*;2QNTJ���TJUD=M֘*V5ñ :a�W���J��!P��$Y���־,�q�t:^nL�/���Mrq��d�
Jt�y�b���$�b9b�W;J�������L^�1Tc��	�q2� 
����OqB䡍+,TK��@b�Ϸ�JȚ2��i�^Ԃ�l\���(����db �=FNT\�+���'
*=�RX�O*�0�af*R�\;��,1h�J�')�:ի]�Y�if+e�% ����ʐ,X*�+�B��[\�@�3�p�Ω[-\*�%�&���J��2zp��{���D�����J$�"K��o����g�s�E��1�;)E'&:eû\�2�˘�R��1AX�J
���� � G���}:�̅ˌ�����.&z\�V���3r{���� �������J�:@C���~��<�M�7���+�` ��� `|��n�ӸS��J)9D�����0%&�J^ ^ŀ*Rdɕ�yH8F��/c �kݺ4 �}�	0 ��:���B^b�������G�R@�TСi�N��%���\T�c�˘�v����B��-RA��؝�1Lb�MJ�aϢ��R\��q�:�����2`7@��Զ�˂��ۥ��Nq���''��ÂDN��u��0@�����Je�]���\��˖�0�壱R��a�Z�wc%�wv������N�qD�
ZX�q���֊ ���H���
w,1DY*�& j�#�Q&@$�8ȥ�\ ��xW4@u%u��0qp�'�K���bıf*T�N*�`�Gsɔ�\�qֱ\�JT����ޙYYW����ܲc�
��&��2lr���4�{� :�LI�y9��a'���{���{�W�ښ! ����h��i�A�HME=E0�ǆ��N������ ��^bM13�+J�J�Jf�2q:���W**U�γ&����8��;ܸ�#�hc�4!�:�<Y�.\ \����2r����X��a�LAD�4�z�`%�
]�`!�dYq�ҮJMp�ˈ%J�+�)�+OK#R�Q6+R��&$	�=�O��FT$ ��J�.OR\d�L�01��u �$&�2{�C]NpZ���2�
�2���eC���C�K�&�0q�\8�.;,�k��R�-��;���.�x̶AED�U$��!I��ػvT�'v)�����@���J�/Nv=1i�&/��⋋�U�+
/A��!A�� ;�ͨ�$0�t��;v1�dÖréZ�2�+��\�2e)R�\�b�@B�����1 C��e�6d'�p��""��f�o�X���I�44�9�AZ�L�#Mѧ8��5��)xs����>]
_��G�'I���:
�(<ԃ9�n��
���X�\M��e.�D�K&&8��]D������t���`Ø�'\UP\!²t��:3��Q�d���sq�Aag�ԡ��R�JsP�N��dF;T-Z�J���H'�*�d:䷸��u"��Z�l A=pH�S����2`
�n�Ԩ���uQ�	K�]mװ3��|@n�E�4b�P��E@GP����C& ���J�d�d�iWc�L�r�ؖ1R�v��b�0ab�ݻ�v:թ�lFJ��uj�ˈ*(� ��rp���]�� !����b�&�k�/! �Gl.�;��|D�*�ʂ�ۜ$��9��C}?����Z�r�+Gv�۷nݻXv)��&���=8��C�� �T@%�3���{����b�,�`oCJe���������B�[Z^W�����T��'�.�e�C��9���s��\�/��P'����Q*�2U @� ��Q�L�*�|���S�є��⫝�v���A�¦LM]֢�.C:^&��P8 � �q��1ݮ{�9�i���%yaخ]p��/�T�\틱��b�v,F#Ak��2Wc��úX��Q ��
�~���Q :Ş���UğϐE�����;2F^2^1'b�P�X���S$2�£(���t��OZ�P�gN�J��#.Χ'�J�q�v��bÎ8�8�8�ݻv���e�]�:����S#!�bt��jX�/+\�daTf²�W#'���,2:rQB�d����w�q�q� �U��J��K��A)7@�7lFv�۲��v�۷n��d�I�Jt�2+9��ΧX��9�4�}	9�F���o6�0�C���5��,�}��D��F���͸.	�f*|_�v���#4�4��-NN��%eU��EgmGVIu�� �{=�CA�������ɦTV
@����JJ��)N/OJ��Z�2�#��K�{���Y 	q����w�w�{���b�e��,Ĩ�A��G3Rr�хWb��vY���e��E�Xb�'T�ZY*�j��B�&� k�9��11Wu�
.�\^����q�>��u:A�Ӌ����8�bg���8\�)iTd���-:��U#�bE��\�<�jR�)ʆL��&M*�۴�J�ZYj��v�۵�X�wn�&\��a�gwl
'F.Z�0�P�KS:�p�1�.\�*�yY�GT^�I��a'k�.,�(�P�t�/#)T�Eï� `1`��/��3�ꠘ�S$��;v�۷e�,X�bņ�d�J�L�J��TC�_��7����\� ��>�O��#u�\�~��$�I��sv��S�Ts��B����L~?��� �.��9P����u("*���L�BA���6����3�(��c��C��R�'(�%,9QD	�R�{gS)2	>�jE�Q	:�$%%R���{���^fLx��c5ҡJ�L���իW%&+;b���ԇ��2*�rŝ��LL���ET�*us����[b�z�L`��  뤸1���`2 d�&�$ �Qv���{��F�f���p�aeBT�������c����P8�<�p�����G�RA�)U�X�3�۷e�1r�#�,2���݌�'#Z�rԬF1�:bdT`����Vذk8�2���X��`�˘8��7S����	`8O��a7� k���X�� �R(QryK�1bŊ�ŋ,X�bŋ�r��R�:�I��5�$�a2�a!b��H̑�	D%Ί��u?�%'������1�9�m ��$9�NN,+*͋�ON�ؓ�Y��u��D�
��-m�,�.��7�iy�Ԓ�+�gd�[�:�d�JS��
`CQ&��p����CT
(��A��Ԙ��NL��Sw���2��Yj|����Zb@���B8���S;Xq�\�@�T��䪉Kb=*c�r�į��g@�c�%Eq��J��,�2Ys���8�/ �W��Yƨ���
J�TN
z�~� �I4�L����&d�q�<�F-v�(�Tˇb���jX�b�Xq�}h��ybŋ0aU��:�u�J�ň�S��L�,bB�9EJd�j��%Q�]LN���4ae�R�=2.t���t�.�w�B��u�dT�3�@�#���d��1Z���ŋ,X�bŝ��re)H:�1�I�.7�+�!��h��{?_ n�YqH�p��#��� �}���y>Àop6d��(Z� �Q[Q�MЇ8����xz9A}��[DUZ�[�a��TG����%��Л�H���)a���	S
@����R�`|�JDE��{�y���QTO]��&�ǻ坻2�؝*�h�˔�"Ϡ�iǡ�4���)J�u)�.R�s�I�:QFI�Ύ�B�D���<)7��<(�ɓ�L�p��MM �_���;u������'���ө����o3 ��D(Ĥ�ꎃ,E(��8�O0��� �$�K���
8�R���lR�&�x��>X�ϖ,X�bŋ0�7v,ScJ�1ҩW1b��.�p�+jR�`OR�Rb2X�I��I�QC%%lw1Oy:d��p7�ؑI7X�����۶+]��knݻv�۷n�Z�rd�Աb��S� /pX���ck�ti�z��u���q�0?I��&bo0a7�sE��fr��������9AUeVgeq�� \fm���3���ބ44ހn���PH0@3x^0Gm)s>LۢEcכjK��j��I� �\d�8�P�K& As`A�P�وĨ@U��`b�Wv��k��v�u��r�W]�\��6 �N���\�v��3���]�:����N�*eŗ.Z)� J�%�t��J��И 2{�L!�\r�{�� ]a"��w[��L��D�]P80I�J:�Q�7�H2��WH*'T{��>�ʊ ���+��GG��۲ŋ0`��L���ݖ֩LŌ|���q���*�j�/��P�Ҩ�v(RР���)&���i�����G���{ȸi�� J�		p���& T`�,W-v0c���q�qݻk˓ZY���JR�<$�������O�a!11P����$~Y�ϒAE��D%W$R#��a�e�}��DY)jn�����cBo�����t�^O`�VU��P#@���ڠ�s��!�����hX]bA*RgS
/
��R	�D�\M*Ԫ!& ��Z�#�/C T��%�a�I�:�ŎXrߌZ�gZ[�]�!�����FQv��YqҤְ-�:�3�%:�t�G��glN��.u*.)%u�?L�AM��*1(���:�2���8��t�:�L��� �:�.dz^�{�ONRtY�$H�FO
�v)� ��z�N �Q2T=Q*�2e��b�k��X�Z�q�X��c�9gT�v3\�Y2�������wn똘��I��
 d��8*y3$��ъ�!:��R2`�������@���h;`ps��)J�5���uK�b��իV�Z�k�c�Z�r�F)T.T&��m{	7B_ ����ow"������)s� �Zg�������t+Y��t�S������,H�y��@M�&(hMI-�Њ��kQ�KP�̥���Pt
hE3=:A*Q�\��R�T�:���*ы��J�����`S���]�ŪS�QCQ�[,������n��ŋt��#)K˄FLt��ыS%����bd��1&)�bjX�b����Qw	zzg[� I�,\Y����2�&���x�|����! ����J��U(��Ӄ��\"����`��#�=IT���LN�-\�L`��Sn���OOM� �bt)��]�=Z���+��ԥv�Ihť��ʄ��I�N&��y�ӋJ�1/%\���tX��V�"�c�	�R,�JJ , �&z)D���0�0����]�kɓ�s+��O*<SyӤL��Os�D�.0�p��bo�7ӭ��}��Z��Mj�Ї�	���8&ȭ��«R�8ۉa�>��j��WA<ii|�����/�A!Ǡ�G#v�b�w���f��x����]'2VO.b��Ur奖�2R���Ԋv�+4�W-.����QTQ t������K�����̘aX��ż`�X�3�Rt�q+� ����bk��ʊ(��F˓;�)�Mr㹈�LK&9�AI���=�^BHϢ
  �&l���:Q�����\́���u��B���%u�A[��T��7eELA��$�*:�a(iJ��&w��h�R)+��S�T�LL��73�wlb�у��:L�T�p���QFCF�Pd��-d���+�
.u�B�K����=u��:
*E%N./K�d�W-v[v���T�*�)��.`
�J�u��  ��u%:0r�'�;��Y����x�`6�"�t �(9�PU՛U]A&�n`��:��*�-�	�gUzDi}�_!`g��S*�8�K�X�	���e�W`{��F�_��&ED)6IS&iQԐ usŔE�ӓ�-`QOT�U���d���kI����p !��X�ݭZ�*�AJQNԓ�\b������Y2R�+S.J(��B�R����)rc�R�= Vy���!����<��盈���x=zs��8ş'碐�q ���@�eG[��q Иs��V�
bz]Z�uإ@ ��Qc�E7zTeE+Kn�t)ծֱ�Rt�f,X�3钭ZTȨ�v']�-������ʊ"��FFN:�)�
�5���b�ŁQ9�8L�Y?5*y�Q� /��rgk��ONc,���c�:ի]�b�k%R������S�(�O}<�a���e�΁������u�$���n��QR\$�h_Vlz7BlPPBq2�<��\/��J�@�ʪɫ;cc��}��ܝo����5��CC$}��U�ăNs6�w��g��H��gTN` AE=*�q�T�JX�:�3+�N A����S�&��ё�v��K��У\^.�{�c���ݖ�,1ja����P��i��촲T��'Z�J��W)+J�@���TS%2JJ��d���.Q`{�]�0���F�7S[�R� �i~����.`�F!&.�g�#�ĹƢM*�F!��K�%&L��Uӂ���X|a4�*(�I�J�2aة,���a��c�L	���),0u��vX��a�X�RddL�!de�N�R8�H:�\L���.N.=1bYj�1�
�	� �R�0�QLK-L��a֮R�+��X�b��5�B�`O*�{���^$��t:��J�Oq�:D@ۣm��
`K'*΀GY���&m��vstU�;啭�!��|�\ϣ����ua�B4nH̩(���g���K�H!�4�m)TO&���z$	%j_3Pt���_댐�ΕNN:��d�u92d˘�b�1ҥB��bĨ�ʮ�-�)Nq����A��B��>�O7��9o��ݮL�2�ŗ)[2q�*)--Z)���GL�q��Z�Q֜X被� ��U-�p�?C�_Χ�����GW6rJ�\ rR�&�$.%g}�	ت#.F	p�������a%�N�)l�f%�����vLI��2�UM�)s�II�L�v)��#��qʪ%ԩ����agcKv=22�J��V�8��T�`��ŤX�:@�T�Ԙ��*L+ HZc�d�%*���T�&T��V�:��X�JL*R	����09��t�4 �0F1	u����6��� =��<<,�����4$�<<�E��Be*@h�dw��ʪ�(��7^�̯�"@ S!����������������R��H��d��(+W�qR�R�rd˗J��T��&*t�V6%��)�'��̡��E�q���c�-�֓-���0�6�U9Hū�b�r�œ
�:z���TŘ�?��(���{��1iy94���*��ۨ�(\I�� �t!����D���@�q�	���.Ƶ�Mr3 ���8�a�L��X
T ��=Zļ�byxQOqe%�):T�˷nֱhQt������u˝��v�RZdŒ� �'��˘�ݭ��C�㘺�U^�)X�c�<��^�i��R�ї-vX���R�R�Jdɖ�L�rc�)&������9���ha��w��LM��.Q{�+�W��� ��fv� ��u����!�T��bGٛb����}��i|��A�Q�՝.������)y:��d��&�7�rs����p���`'�B���Ұ�T��I�11`&T�T�R�*���ˎ� ��je˓1��!%t��J�%*H�`w,3���*����Qp73�=H����:�ŗ:���ؐ�*�U�&@C�~�Djt���6����3�HDD�8@H��f\�T1/}�*{�#' t?��D��KK2,@�D8!��^����EDeC 7�00�Rd�l�R��X�`N*t}ib�X�R)J���-JA0�H-�1j�jE�2P����˘�w��H�s�t�Uî
��+ QK�X
�(8t��M,���0`��;�d�J�L�J��°%&))R�� ���z�t�@�OA�e�/�����t�ڙ[�[PM��&�Kc��M��	�A��Rf�x_t�JM�n��EG�����}��]-�6���a�q1��ӌ0H18I���^�4BhVYrO\A9*�j��D�j�I�*)�)�)�) AH�.ֻvŉa�v2YJ�`���k���@	���|g�jI��J���b�0#CC��.J�0aV#�&İ�]�R����5)�_�X�F=N%p� �t�����$���!Q�l⧮�q#cGڠ��rQd�S��U�D@�*��	�ú��g9z2�����&MȁU3�b�� �8��J���v�10��喖��zb�7q��"���R�UDc�S�q�=JX������Q���kTL��0!�R�]�����]�;,Xu˘��bɔ�J��b�
�*8U1���n2W�I+����<=�B.s5���侐�D���nwQ  A����Fy>_�
���'�B��`͠�D5��	���R�$��jIzYy(8OCR^�JY_�����Wj/�1J��*#*�J���L)� S�\d#&T�r2yU�T�O`R촳�Ŭ]�Xr��ˑ��ZA��&@+����Г�,3��L�D�6?:Z�,��� bb�a]ݮZ�L��du�V��TbX%���� �T������ {��/�u׺20Pa#G���0�Д����Ǣ�V ��bON4�*&�Ju8�9J��s��J�taKR�L.@��{�똦b2�ܴb��b�E[��r��`�Ԗ�O
��ZYqf6,X�bŋnݻv�۹ԣ#vt0�q+^U8)���TRbŋ,:�+X�\�u����(�aK���T\Mi0�&Q�绝U���jhzs�:^Nw0�R�ZK�)�Y���]��}	@�b�H����f�y�=�MBO��%s����0'�:Kk�Ϊ�n�!$���/�52�9$�B
A�Ow�����DW@H|�3����8��e��'0
/2Q
(�����`�ybŋ,X�0`�ŋ&J�:�q�*V3�X����E~�`*�Da1�̘�����$�F]�u���
���[-J�O)P�թI���ݰ ��ˊ����������PY|�CQ ���-�%PҐUCQ=9�KєPª'�>L� �]n7vU-�@M�J�)Q��s��	��FJ����;Z�3�wv�s�k�Yq�%��a�Fn�r�S.Z�rT���FRX�2s�l	��Z�jիV�,X�bŋR�@�R�u�J�)�eS;**Ě])6%�,�v+��&���c�LT�����8�	��+:A��^�-F`N�zK+���3Pq�<��ϖt%b�sK(3���q�C�\%��t�PW�[��T�H6��f�f�y�9�O�SKJ�cc+�ue%]���}9ƀ��'���R�_zn�D�D���<�t�YR���&���L�U)�.L��T��K,X�bŋc,X����
  ®�η���c ��Y���t���c�]��,�ɥ�ED���1�_���I�:��T�1|ȭ��= 0.t
9�((�>��XU�H0V�P*"����z�eD��	�����=w�Q J �3q�)&\�1�/,(�����H�.Q/b0���K&L=2�*�e�G�-���F]��;���lI��Jq�k��L���v�۷nݻ0`��TQ(��W�� rT�����R�\�we�v;�I�*�r�,S&L�f,J�\)8�s�W�3��&�|���a� O�G�KcQK����D�!���$0�9��u=���a�`O�h�ͭ�"�a&�B@���V�����ȋʯFnev�Ԗ�S�Y�$�6W)Pq���p�$�d@����	u9���JMP���H'�*)Jt�өT� ���M2�ŋ,X�l`�����G����a��w��?cF{=��7Z_��u�D�%/�ZM�&4 �\���k�կ043D⩖�:q�zZW��H�CCt�:_.#׸�3G1eF{ �R��Y=
H�,d�rps�9��m6y���J�LA�J�	R�%Hp� S��s�Ү؆U�ݝ:�ĀV �F,[�LUie��1h��l��;JRkV�&���9�`��3���X��3���)8���w�|u��,Y��+�b�*S�¥:LP�gR�v0�yх���
~�u?� �(b�1Xj����e�}��Y|����fE��d� fJP���F����6��VUg#5��P3���.�ol@W56rt�@B_@o�`[��ݩ��q����G;��4�ir�?��gS�*L*rs U)I�`
@��b��*����0f0`�ŋ.�F' >�ouu�x���~đ�_v�f�.�5O:^J��9�Q�:�#�	�M{��Ӊ�Ju*S��B㋽��K�gN����&d؈:���$����������!��ˌ@��K��+:�K��LB��LD�I�B�T/`JA9Q��N �Fs;ʩ1%R�P���rѕ�T�v:p "2d��x铗c�,��c��G�L��q�%��U��ҫ��딖v�b�L�֨��Ě�q���-۷c�\�`�W.Lt�S��&u)��W�TE:�FHn�7Ӎ��{	�9�E��'���W�X���Y�z�3/&JJ�X��d�����a�u��gI_Y_XkEa004t�QQ/�:#cS���y	����2�;���i~�� �rr�>���V���X� �d��u3�H
 L��'J�R�q�0`�`���c� #���[̹ކTQ�K��c�p唥Lu	�]�t�.[���Z�����,R�R���QgQ(PbXP���r ��C���\&�a#)����XD�XqB���c�b!Q�QNZ�$$=2�	X��9��r3F11TFN=$t�\YN9gki�-RAH�����Ö�b�ǌ,�bս�d�5ɋc��\@��b��[���J�Hs��H�� �y\���0`��v�v+�.R�p坎�2�*T�\t*��A�,H� |���>�����n��t�Y��t����n��`��X��r��4!��)HoiYP{2� ="�B��FtS�2K:J�{�ѱ�!��s�(,�#�)g@���))gS��\�&��V|���R)QRU�J�(P�X�L�r�c0`����-�w�.΄�=���)MLƘUjձ��FQΣ#
s���:�R�`��R��1Z��y�b�J�,�)�š_�СS��?��L�Eß�Np3��	�s���0 ��~�)Lz.{T~�T%=q�=<�^���щ@_�a��h�ՓƅT�H��B{�a��9����Z(-������,4�FT�w�;v���ҧv+~Yjb�
��\1m2�����0a6*I�OO J1(�t�	t�ؖ0q�,8�����R�L8���&L�2dɒ�C	 z&M��$������dz�s���_@/6�g8k���/1{���o��ۜE�	��f�t�+ �q���&���1�c�����*���h
�ntCƅ�KCb�8�c�kK*��;	�K�i��!�HM��bV&�SLM9<)B�@���X�\�h����-,8�bZ��zi�%�]�Z@�i���_���Iq�b��T_O2��V��T	�1R�K�c�X�.�!i2�;L �2y?�_a����0aI�+�}�Q	C\�O"- �04d���45�fuB��&�p'�	�@b��֢ �y� �:CA�M�otu�����%)�E
JT�b�+J�8��d�q�*1`����-���J�MZ�{��aw��0]���e���0`��X�NQTFS*v��[��C+v�af,Kv8㎵�e,W)L�k�N�:t�ө�W�ٕi�����HH�n��^N�A��4�%��`NT d"�JA���eiDV3$xIIt�3��59�D�]��#���PDGHWxYz9Hg~��MZFk@N��҂�(����B�K�:!#��Y>1j��0U�I�:MD�*f#��r��W.\���`������0��)�@�B��&�Zw\�|�e�j�ʡ���\�=F~��	cփ���
*S%OL:�
k�Ԗv�c�G�� �K�@�Hq4;���u�:P�N5���J&�68_�D�шTO��'!� ?�nb����1����q��`iIJ�K���~����ba���J�0��%%y�S��n�uǤ����W;��Z)��d�I
V���a��񅔏�,���W�z0� ���˕N�'���v��b�J�R�%2ի��`
L���TbRuK�]̒�B@}>�J-ɲJ+`k�RQD֓&dU0��c�	�.�n��/":�]O�6�;t4M��Rf�4�l5^G46GX6_s+6/�2�����"�	�6�7W�� �J^�O� w�����%�xJs��f%B�J�rVi�,Xv!N�:��0`���,0`��b�)��1��J�Bu+ܼ��2rf�I���>Oj�c
�ZF��kv*T@BBJ%��X����-���Y�~��[@�OJ���V{���N�ˏ]@N2��C�qt?�!�E��L������X�0���e3{*8��NW�O��K�M�f�u���'*dJ �tG&�, ^��ԧ!���Z�+`���OW=J�=M�S\(���g�#�h��K���d�U)2Te%��:�uɹe�G,1��+X�*AJ�(ĦGV�Lt�gV�.C%:�,L�$X)p����_n�/���	�=�+b�|��8@�Bd���s� #����I@s��<�����J+&m�A�j��B
#ɺ�ms�� ܖV[�1'�GC���Q=y*�9��ѝ� us���˘�Z�j���
�����0aa�0`˲Ê��3����:�(S"�����t�݌{9(:��* J�.O㗈�� �Pݦ`bM(����uh�b�Χ#�]8H��l��{�y�����A]`�bo0��#���t?���w�T4�`�q���!��4e|�#��E�	@�'���v��0����q���:ğOg�aTP�IEX�*���M2ժJ�-0g��B���F]���3�=N�dz�M��2�R�)��،�vXc�)�-�\�3+���R,�N:T�P���R������CC&z�T :��3/_|�'?�_�p�O����v�8��|!�f�ʠ�x�Ĝ�'�&��6sU�5t�Cp�f���Yp�8\+��M�CK��e�&���Q��X���m}	�/5�>�o�7�ө�� �ݏ�\�Jd�Kt����3�0`��0`���R�Y*{���H�2u:BEĝo�*rrry�#��UXE�@��n�;�ɺ�bz�}	�˓& :�ڒ��'���a/�'t�E����%�"H�q���A�n������:�@@���`�g�ä5�$�X{:�b��Ǹ+���8%����Ny�'��[\�.��T� U�rdɓ&L����T�����,1N:�.����݌�N�:\�t�# ���Å���-R�.UM*U�V�\�wlS&b���N�T.FOF22Q`
)8zp1HC�S��Y���� 	y��\�o#�0 `g!0G�+�Ȥ�\i�$"H$"H�U.	�	7A�n�f�(А��AJI�B��ɺ��}��\��
��p"Qv�`����������
,UA����|�46 �R[;���C ��hť��0`��0`����v�t�k��� }��7BB^�﷐C��H&�t	��A�@F��ʐmt<��].��k�5�&A1��)��&�v�C�GZ���C	Xs���F` Fo�G�k�� H8��d�CQ1	.`$u:����A�߯�4A'�)�������hβ�= s2�ʊ21�� C �@����ˋK�,[�l`��ņ�qj�e�a֏���;v[v�JT�a *"�"E����v3�V���=�	�\ň唩L���$ԅOT��
&F(j!H
*()��h�H�r�0�WI#k���A@e|�8�^A��e;�0@��^�Vzj���<8C_`�Ī.⟠��H�&k�H�)*��ogC�$h��A�f&�U<j2`YW�Gp��<(���gXOJ H		
�q�eW;�,;�kT�Q2.N\��b�?�0���0eiggT�@880@� $$,�u�Ĝ��/�`��؆>U%������/!�! ��Yq0�ꊉ����Sc3D2��0ti`�Y�&�{=˝"�� ر���5���\��1����H:d�D���d��;��z�s 0:�d���ә���2�lr��v8�R�*�q�Ö�,X`��ik���]�`���,2Y1���ᇯ���U'S����JL�z�1������Z��T�G\M99E8�2iG ���AJ���o���G�W[���� �Bnܞ[�vŗHӄY��XYt��6�ޚ_%--��u��b"!��K+�YI��a�wR���@��˂���rGD_@lPPs	>��䎂G�5����bd�f�xVUs >�BB����ϗ��<�a�%&L�R�W1LM9P���T��Z;��?0aa�0`��2��g��7K���OC��O7�bqa������4	�&��:�\b���c�+Gb��y�s+FLzapAuC֠�טs�� ,�y�/QTN "�Qq����	����0�E.` ��AwY)p�U)KŌL_����/ь�����y��������j*��P��a�ǌ\�2�J)�c�[�,X�a�4�Ìc-������w�JLY�J��+d��U��d�U� �)T�X�R�r��T��9��1EX���u��A��C���ၣO�+����̀�����r���=$) }�2
_o7�t��ɩA|5�⪾�`ذ�j)q�=��%,�Œ9��Y�՚^������NY��Ɩ@�nv�V�0��c�=��l�_)IXju����E- �%V�:b,dLQ3�R�*M0�R�L8�1Z�ό0���0d��n�q0��$��a1�0!43�E��X�S��
�c��M.�z�q�%�[2�c�\t)z��I�J��"�H�&f�V=��C1s��_`**�!H*:�K֨��:�(�'0`z)	. ��0Et�95I�z�'N�{�=�O07A�zy�z��z��(�����]�i�,[vu�bņ[2�0w~�iaح-��w��u=®T{	.C~������R�p�\�)8�U+G\t�7k�� @+ ��)RLRP���S)&�u=ʺ��e��.��BĠ���[��| �iY�	�A�.R��y��#�P.aS���ư���hx�f�IW9Yt��\���P������ʄ��h��}��N�0��'
   �SQ�������|�>�O2GS�}����|�Z���E�� L�e��&v;֦R�s݌�,0`��Y���X��R�T�?���gH�>[Z�,����u2���]�T��[,S�0Rd��`s��$ ���:,�&4��t=�`"�iH ��������` �Ee�,@S�����&\�r�eK��/�A@��j&)��O��
�Q.:�)p�X�v촲�ɓ0`��,0`���0`���0`���,X�a����	T���B�6�#<�n��_�JK��y�+�a�qU+V�Jt��S%*@�Ί*��T�gG�������q�/)ms�Z� ϧ�5���f��&�}�_ ON��`%��2�`i�YB.	I B�AI�c���6��s�7B�M��CNe��U�0)�eͺ�X]��q�?�\-E mF��'0���u����s>�՛�Օ��D=rZ�JT�IW-Z�3�G���L�ql}��뵣��F,X���lX�b�+���`\2[�--C{:��㩟�N�у0`��0`������F�cF	�I��A+#B ,��70�{������&�Tq�U�e1rP�TQ� Ę0*��X%:X�3�������Q,�)hTɎ�1=��E:Z���cŋ�0`��0`�����,X�a��I����Ld^�U<$ �� �8�e���
Ā�f�zs�*f.�b�2�ɔ�:u*���buuh�Ӥ���LT��*=9�ԕ��c�|��$d���rz04p�"8#h��H�h������J	�h����izz<d0��L�g�@�@�/�c �Ck�̂�Ԑ�n��s�4��5$�?P<qr{9�j)�_��A�	����|������*��()�X�b�*R��O ?v�r����n֎[X�b�7kV��r�� "��X���>����4hiQJx3�i�0`��0`����,�I�:�FSF�lh)eajp��I���Oי��@�Q�UL�_%���yQB,�':����P� �7d��P�-QIaZ9p������{�Ի:��KcÖ,�q�0`��0`����X�b�%�,X�b�.�'����'!��L�\AhP�����J�"Ɋ�s+��L�JT�T�b��5+��	T�l/�J�����)�zb�}8�O�����g[���	����R�Ճ^o�g��L@0�X	���{+�����#��/���A��-��vt���=t�ZJLLܞ�F����
���4�8ɥ1J�y2��+���( �^`��W&RM��T�V�L�*T�T�MQ �1R
G3wv�r���ŋ�wn֮�` ��a��� ��Φq�ۤ��e���Ɍ0`��0`��.]R��`u�ҹxC��UJ��lB���L.H"�Pzt�� � ���	Sԋ�:C�¨�8Ʌ�����������Q� �:�z����`��	Q��,0�����&J���a���0`��~0���0g��abŋ�v�۷nݱL�^�u��
���	�:��D��S\12Qg3�*�#
�Rt�QET�R�*��X� ��2�\��c�R����$����/7��uɡ�@� LY����/Z�I@Yms�9���F&Rb�����A�[^[M@�MA�M�����u��3_Wd2���O�E*�Nw�3��� �d5� A��}��@@M!��!��7�(��!�rz=j�$Ω\�k'T��)&bM)I�-v0gݭ�20�bņc�1��$©-�]�*Ł�� �u���T���0`��0`��Zt�f+R��+ ֗@T�B���1;�H^TLͥ��MDS��T����,z ��{#?�/%�TC��qaOwk�B,��\��bA<�V5.�E'J���0`���v8��0g��abŋ�v�۷nݦLT����ňJ�t����TR�
(e��Β�J�1*S��*�re)N�J�K60��I�'Fy�D���IN���<�,,+�(7J[�sFCK���e54_a)WHrYjQq�_���"�1��Uv����Ҫ�#b�庪�R��q���U����PPM�\G
B�+���@Ԏ=����\�J� �鈂#S����R��Ҡ�.UtQ�X�v��2i�;\^(r˒��b8ϻZ9ldabŋ�-�vU�*��rŝ��yp�X�)l`��0`��3�L�4bXǸaR�A��������),�_���q�����ӃOH���2z�)`���MYƨ�ĔX�=�0���y�]�QZYp�3"lV��v8�W)\8�f0`��X���8��0g���0dabŋ�v�۷n���LS�C����Z2�as"
k��`��q 1b�W%L�r��T�R��2	�:�z,�1L�\�~��?�с�i�AÇ.p�=5�"�2� � 2���Nw�tv��3t�����y����>����A�P�^W�[ܚ\F���'ua�|5���X�\�~_glXB9U|����#�3���o"7��>D_@�!Sv�0����֥sƁ��Ӑ�V)N� T��GH��R���.��钦3v�r���ŋ�v[�Z�(��X`�0��ݱ2u���R� �[0`��0`��b��*�f6:��P�S�E���*�ڕB�)2G�1�萔�8�]�)�2ɔ��)�$��r{��?�	��L��-b�i�0����>Y�nXgv�r��f0`��3�v0`���X�bŋ-X�b�%�,X�b�ԓFy�.$s<����lN���ړ�`������X`�U�X�J�H�AB�L� �R૖�*\�~�¥.`Nt�<#����JTO��d"�+/�#ǆ鹻H,m��xxYu�'�=�L�D��B���#��ڈn�Ծ�R�PW0���R[ЕTF�%���j��E� ���O}�+�C5e���A�:�*�:�	��$�p� �56�-,T*��J�:�)4�X�v��<�U*W-J@�k�۵���F,X�̳�ܴq�]���k2����% q��0`��0`��KaV�u��UEFt�ɺ��Ow�K��D��bz���1$F)
��de�J�U�� �,��%�$�� LV2b]`
��jR���GF=N:��X�3��q�#0`���0`���v�۷n��,X��bŋ,X�)q��8�U�gC�92z����1Ϊ>�B`B⑋H\�IRd�TTS�J)qQ`��~�'�?C�\��l�)  F��$f�hx�h�t�!	�I^O�"�7Hkɵ�dm��q�<�Џ�^ ��ANg��ɺ��B���#��DT���P$s9�\�A�Й������Fg�x���QV*�G@�ߣ@ �g t�KV�RT��ACR�F
�p��֮JL�Х]�w�Z9ldabŋ�v;�Xbգ#>���i�@���� O!!d��#0`��0`���Ի���:�r��� ��Yr��G�K���{�:��`$��#u�RtQT��EJ�.�@�e�wk���TKw���.u�#bZ0*ԣF ���Z�g��0gw:�c���ls��u�zh�X֦�%~�IN�b�Y*g������-�<�ì�����IS�S*t�T�R�OQN`NN` t�d�J�)P+��� :���.^�h���W���A��DAXeGDd q��Z�p�^`+��
�O�֥pZ"*ʀj�S�K���y����x�6<,!9���`��1���&\�{*��,��$:���L�Vu�%$~�8N�@=�!���"M�����)��`
9�����.b�rdɝ�v�J�cÌ�0`��0`��,0`�`��18]Lbe��]��`��1vYk�kwi��0@�L��g�T�α$��W[� X̎����U.Jt�D��a�WQ���@ g���LS���.Q&���1Uɔ�;d�#���;��?�����n�
ZZ2�rŹb���!J�!�-�w	=�Ɋ%`JA���ɓ��- e�J�RT�gJ� L�ӥE'�(�-�թ������aLB^a$���������m@�v���͚��4=�g�c���	�:�QM�����
�rC!c��C����lxQ(CI�.�R��;� ��!%����p�E����BaL��D�d�'�L���((���E��oh1F=t>�]� L�DҮ� (�4�%˘�Z�r��-�s�֭v30`��0`��,X���1�0`˵ܴf1�o�`��1j���;ߝ��?Q�� ���H�Q8��� ������b/u*S-v�u�j�GL�:R�OI������C���2 �$�QӢ��1:�+���S;�-����d)oZ0��c��(x�Ә�w��K\��kR�1 �qT�X�20H!�C��a��M14���L����AH)3�FK;v��[�)3�@'�)� ��XD�RR�VPhk<~�8\�BM�7S��&&�q�������v��W3u�e��i}?V��N��)�]�R���n�8��B Ď�0�r�s�ͭ$��Li���묵+�J�q9׆����|�/ @�:�cC4�"�{4��N*�I�eXɅO�14�˘�Z�r嫗�f;q�0`��0`�ŋ30`���c�J9l��c?�0`����Gb�ṕs���֝NR�`�	�JJ&�o��Y\�A4�Ԯ�J�X�r�Su�!��/t2,S�����u����E�H;Z�,�jeÕ,0��b���g�v�je)��;vXv#�)g^���K-dQ�haL�	� M3���q�IB�./=�?A���ڞ"������R�JT����H MKiR�:�� `kؕE�"�4bH�4��������
��G�i� �J+���jz)V|�!�L۪ ��7ɛ��l�]̊�ek)V3|���F��SG��sF��W;��2��B#(��A@L!��C�d��@X�ٰS���@֢��ѐ��n�<�7\�(�--N��íL��ԩ��d�&ur�˗.\�JS�WĪqU��KF0`��0`��,0`�`��0wy7����T|c��0`���-�7�(�)ԙ1L��_�O2�ΐ�gA���R1x�J��#�- N12��GL��{��
R��D�d�u<�/�'��*s%��ŅC�ݭ���0�n3,��Wq֖���V��)ܪq6+]ҕ%
��u�:�o��%����F}b���\� s����S;JKœ����H�ɓ��b�%:��~�:�J���@F��/
���OK,�T#��һI�����M��lW_l@|V�P��/��"�t!A��leja0h|���J"*;Y�+S+AIɘ�Iю�O�Ѡ׆P7Ypr��������D%���1�{��5L��1&�h�s9��e/r�!�7k�Ԥ	�LtRf,J�'�bt�U*R�:M*d�I�L�Lrû�0`��0`��,0`�`��1�:z+�c���0`���L20`����% �j�$ҭ2Cv&�bd�.%	CL�I�^�a(ic���`���)1A���r����b�̀@H'����!����1et�����ʻ�w���Xq�~Xq����F)�D�K]�=FL9jhIH{�Е��$0���H�id�K��D��'Y4�)���I�eH&t���ԩJ�M*d�I�\U%$�Uɥ�DI���W4xG?,/��͐NV� �K��H�f����x��&�zjmU<U4$V@Y}6�8^������ʈ~@xrs>�`�AA�������|�L�B�
�ƀbJB�8�	�$�������ƅ4+��G �H`�UWJ�}����Ur�%V�&UIU�R�J��R��Z�(��]�Ru2у0`��0`�ŋ30`��b�c�+F}���0`����K1l`婉�bXu���n�"�L�FN%21lhy�?�M��	T�۵� �{�!cW8�qz{�U����E��IE���+" �!K.�J�떌���c�,]�ػ�8�P��=t
�bP�(jK-� z�^J��dJ��J"f��bsХΐ7Ax`rRi��RU(T�%R�O.{��� @�T�S.L�1R�G;��݅��Y�b���l�U3<"5��������^l"�U���֡�8ә����Vs: �&�*$ !�ǐ0@#��y6됊)���i�}�Y�L�E�z.�mz3 .�?�I^�/1s��C���㔐�����y�]Nf�WȘCuAe�@�YAo|���A��T�LT��3$�.�'��R�2d�R�:�r�<u$
0`��0`��X�a�c0`��j��,�g�`��2TQk���jљ5��ç'��%�!-�>ʎ����LZ틲�⒧0'���<������A��E� �2���Ꭷ�SЕ���\O,���;�����3�v;����O_��^�E.Z���r�1ԫ��8�O�p��`��gS���A�a�!qwИ23�ԆT��+��F/d�z�F,�JR��
U*R��1��&��s�8B�H��H��	�g_A#3F�c�
����aV<s�OMVڞ�_�CBo�� 5�W�G����q��̾��F"5��_*�w�ĖB�Q� ����9!��)��9YP�����U)346XWaA5	q�
O*"�&d�� ��!�TOJA*c��.�\�j�+�00[�.:()5,X�0`��0`��,X`����0bђ�U��w�0`����{0]��\8̲۷qҏvT��/��z�1�E�g����Q�Ζv�L�Z�Qr�K���t���&Z4�q���*S��P�E���J�XuǪ���0`���n��we�c�Z[���Q�.�	U�kS1-Ҧ� �.d.z��Ү� ^�	\A��t8�E�������B����&E9H�b����� ��P��I�K+�iܢ���{��RZ��Z϶�}����.s 46�:]%+-���%�2����s5��?\-
�%%.NqǙy���!�r���AH���5q�Q�Wp�l�117�I�� f��y"#��MO�N4 �<�Zo�sƐ������/���l�9�%��bM8��d��:���T똩�q�u�S)R�0��}p�f0`��0`��X`����t!���e�,X�b�ݖ1�"���e�K� � �\�;Vy�FkS/&�������p��a$�X E���x@t��1F.J���U#�Ê*��0`��Xq݌�0g�.Կ�	�]Ou�ɰ-��-L1�*� 2G�;�苤h��y>�/s��:� a�X�vA�=1f$�B�b���jJ�
QB����?'�v�8�k ��"��|�<��׈�٫(�ͺR��	s����� A ��g��
��k+R���!��z ؒ�^4�}	���j��%f�������+���� �V=p��o'��Ɔ\4h��t�7�0�'[�����jE�uf��#��5ea0d����1E@X��Y���dĩQݮ&A2b��L�q5��S�S-R�X�gnݖ���0d`��0`��0���?��c)�W{�n��X�bŋ,;���
�b��f)�TT�Q+��X�1�,,�'i�Z�2biN�10�:,,Ɨ:CD�O`X	�F�gn�{��0`��;q���L2��d�H��/�ᕩ��;,2Yj�����L�o�І�� vVǱ+��(�{�E�f��$N�-i5�T�Q&�u"����`�IP�!TK�m&c�"	����mA<���P_XG<mDn�&W;R�HC���u�49���Z���]-��Kܑ�e�x��Uh(�����L�����u5"���N�$G�I(�,�M�6����t?_�.`׻�| ��` ���X!�&��@e{4�4��=/����>Z_ϥ'�v�JU�E-J\,�(QV.Ҙ�.L���ۿ�*uKc#�,3[�0`��0`��,0`���ZY22cXq�K,X�bŇvY�鎓	2`�[�B�[�u=����,ab���҅FQ,�<���%:��x8!U�b�̉_��A�S�-v�fY�����0`��v��a�?Y۶.��x�����]�Z0u�T�:�p��HD�E�H^�s�,��* ���S(�B ��(�f�S��A2�*H'��:���)rԢ�'9,,,"��/�/����L�*�
�-�����k'�G�!T�^��O�]��De3iy>_��f��1fB
�;�
(�$ZBI��a�˝�!E��1s���"���q��Q������|�����`������a�����H�FrUt:]E.L�`�-���ǯ�#6�����O\:���R���
AK����V�L�1Ja�R��<(QD�b;��v:ծ�����0`��0aa���l�2yT��X�bŋ,;�ŝ��pW�����qOҐC ]&K��TTS���bđ� $���=H �zT��3�d4ߖv���c?X���0`���,�u�F���=D0*����vŌQT�H*�=�"��K��U洕�M��u��:�.��&SCEw[���&Z:bkJ��(�L()�WOO:d�s��*�9ՕV\�*�wP��:*J#��]Y�䈂����h� �)lr#�#8_Nq'ӑ�8���Ύ� �`�f�frp��Q��������n�4��狔��_>lRЈ��jlV|���:�ߧ�q�`���h;���z��\�3s<�n7AR`"j�H'�N2b1h�)(�el]�L�2�jR�vu)baX�ZZ����e2��X�L�*�e��0`��0`��3���0(�1-�,X�bŋv�bŋ;�����0:��X�p3���f"�R��[���N�㣿�ˑ��0=����$�9a��vXg0`��`��3��ݻv8�V����.��Cie�حZ��bU�R�##��@��wCQH
WCuF�^�u:g�G����/`��%,X�LU) �S&R��1B�
;�æ �d�@\	��a��H�UgrP����NQQMVQ�Q\�@���^����q���eT���zhW3jUUlf�V���ښ
 ����KS�[z�3Ҁ�D����`�� ����	������ր���hy�� ��� ���T
].��o����n�4���7ɺ4ֲR_�
��0U�kK-*�)2�VԥQ2*�3���a�0`���1b�2����l`��0`��0���?��:�Jz�#�K,X�bņ,X����+bz)1RE�'Jד���������${�:�u����(�RtPWn�Ê�&�`��ݦ3��0`��q��R8�vX�h���C�ITFc
�1j�W��L(�Y��Pex)zxs�E�A�d:�\�p7�:�"���Y9j��WNORT�d�(��*���Ö\�P�+��Բ��s4��=!����2��CL�\�,����K+�hmH) jˀ�A�6s��DיЕ��
�试w�5+ �U�D�.M�07��X H��� ��_�O��@Z��
9������hh��q$,8^MBb:jT	}�^hn6��0���������4l�PP)4u��(��
uie�H uJ�#�JuPĂS�e�q��jիG۱֮Lu0�ݻ0`��0`��,0`���,1��%T�Rc�,X�bŋc,0b�b��������?̜ĩ�wXq3%�p��d*yT�`���D�eN�CJ@��$�r��X��yb�`�0`��X��æ:@wn���vTA��/vYs)wlKuQ�F/p�3��"u���/{�%}��_O�S�Lњ6�.t\:QDҩOJYh�I���JT��S���ӑ�<��^����ʫ���p������y����0�49+�Ö�\-G��೴���9<��W�TǂE,����l�	-��.p5�����'.M(#jϡ�Q �evP�3A�KR
*c���l�$fh�"hܬ�ZZ�_�a���ꀙ�������1� &�=~�#�=�$��'� B�p��U����)`NJ�)�9dɘ� �3 �lW2Z0��ݖ,0f1��X�0age�0`��0`��0g���Ω�Q@���bŋ,X�lagn�v:�r0��p�ld�A�%E�}�}<�¿�]�:�J��!����"�₩F=/�0���0g���cr��u%��)��V�\�b�Z��jc�]�b;��WY�W��Jıp�� @s ������Pr.�Q� @�2eJ�*��$	�J�2R��̉L��!�=�A�j�bA$�(��D�aH�02��p�g��H,�kkDs�6>�ȩ���ܛ�b̠92�3����\��[LL���������P�[���u49�W�f��E�m!����Rf�jVy�MU�[�h�X��E�������i  ��d���o��W�uY���x�3u����C��&t�{���12e.έ`	T
���kX�c��X�v1۲ŋ0��n�q֎X`���0`��0g���8��RT�ӧ]�q݌X`����,YpT�
W.*(*��)��"ÅC�8���㡗%/%CT1NN	%J���0�	�
]�vX`��3���:e�Ϊ�)Zt*�2ШjS�TI�ON&����T�YjT� �d�ηX�*2��C�E��y���1:�`j"A���@�eAB�
 @�2l��RT*y2�T�JT�$��U?�E��ߡ�, "җ��H1��~���̟ϷC[2hWB7jt��:��!d�'͎���u����8��tI�"���s,M�VR�����j��{���̠9=� �U�MZ�UU[U�[*́��b��ӡ�����)pC��/�����z��,�z�y(=9Ĝ��\b�2�C�# �(�B��
A����b
X�v����;ZŊ�c�,X���v��㎴r�,X`��0���?���v8��R�@��֭�a���,�q�t�U�e��I�)�����?_� '��s���aTR�ߠ*�I�=�K1]�3Ř�0`�����1IT˒�`
�H����;��T*0� �td�#�J�k��ODAR�1TQ*�!@�鴥�$�`V<YUBg`b�(P�E
 A=��2aSщ�J�JR�ԥ
Aq4�g�O��5D�jH��@�ϡ�"������H��J)�;��x��Ԓܔ$}��_nN��&�u`[��$"�|�5�=��2���9Dl���b�f��Qgge$_gXG<9qQM]O	.#�j����\ ����$s>���
�|vX� s��]�z��M��~�s���d
��OC1FN=O2*��N:���kX�c��X�v1۲ŋ0�b�ݎ8�G,0`�ņ0`��3����c���`F`*�k,V�v���v��ū�,�8���ɒ��_NRP���JP