3832
500
355
3
0 0
116 100000000
232 100000001000000
223 100000001000001
207 10000000100001
238 1000000010001000
241 1000000010001001
231 100000001000101
212 10000000100011
234 100000001001000
243 100000001001001
213 10000000100101
216 10000000100110
245 10000000100111
191 10000000101
165 1000000011
15 10000001
20 10000010
147 10000011000
196 100000110010
229 100000110011000
214 100000110011001
218 100000110011010
219 100000110011011
204 1000001100111
156 1000001101
122 100000111
18 10000100
52 100001010
143 10000101100
188 10000101101
160 1000010111
128 1000011000
182 1000011001
55 100001101
117 100001110
118 100001111
53 100010000
175 100010001
21 10001001
115 100010100
108 100010101
189 10001011000
187 10001011001
183 1000101101
56 100010111
22 10001100
23 10001101
174 100011100
101 100011101
114 100011110
57 100011111
184 10010000000
193 100100000010
205 10010000001100
247 100100000011010
209 100100000011011
210 100100000011100
239 1001000000111010
230 1001000000111011
222 100100000011110
217 100100000011111
63 1001000001
65 1001000010
104 1001000011
31 100100010
95 1001000110
136 10010001110
131 10010001111
98 1001001000
179 1001001001
70 1001001010
153 10010010110
133 10010010111
30 100100110
28 100100111
67 1001010000
173 1001010001
68 1001010010
178 1001010011
35 100101010
135 10010101100
152 10010101101
180 1001010111
29 100101100
172 1001011010
105 1001011011
6 10010111
1 10011
54 101000000
111 101000001
177 101000010
112 101000011
4 1010001
24 10100100
103 101001010
123 101001011
97 101001100
62 101001101
60 101001110
100 101001111
145 10101000000
197 101010000010
198 101010000011
192 10101000010
228 101010000110000
242 101010000110001
249 101010000110010
235 101010000110011
246 10101000011010
215 10101000011011
199 101010000111
110 101010001
121 101010010
109 101010011
5 1010101
59 101011000
94 101011001
99 101011010
61 101011011
130 1010111000
154 1010111001
107 101011101
27 10101111
26 10110000
25 10110001
176 101100100
64 101100101
32 10110011
8 1011010
113 101101100
58 101101101
102 101101110
106 101101111
13 10111000
45 101110010
119 101110011
3 1011101
2 101111
33 11000000
34 11000001
7 1100001
72 110001000
92 110001001
137 1100010100
132 1100010101
66 110001011
9 1100011
36 11001000
69 110010010
93 110010011
96 110010100
71 110010101
75 110010110
90 110010111
10 1100110
138 1100111000
134 1100111001
74 110011101
37 11001111
11 1101000
38 11010010
73 110100110
251 1101001110000000
252 11010011100000010
253 110100111000000110
254 1101001110000001110
255 1101001110000001111
233 110100111000001
220 11010011100001
236 110100111000100
240 110100111000101
250 110100111000110
237 110100111000111
202 110100111001
200 110100111010
208 1101001110110
225 11010011101110
227 11010011101111
185 1101001111
91 110101000
76 110101001
39 11010101
77 110101100
83 110101101
40 11010111
89 110110000
81 110110001
79 110110010
82 110110011
80 110110100
124 110110101
46 11011011
43 11011100
42 11011101
126 110111100
84 110111101
48 11011111
139 1110000000
140 1110000001
171 111000001
49 11100001
44 11100010
125 111000110
141 1110001110
149 1110001111
47 11100100
78 111001010
201 111001011000
248 11100101100100
211 11100101100101
221 11100101100110
244 11100101100111
194 11100101101
151 1110010111
12 1110011
168 111010000
186 1110100010
150 1110100011
195 11101001000
203 111010010010
206 1110100100110
224 11101001001110
226 11101001001111
144 1110100101
167 111010011
14 1110101
41 11101100
50 11101101
162 111011100
85 111011101
169 111011110
181 111011111
146 1111000000
148 1111000001
166 111100001
158 111100010
190 1111000110
142 1111000111
16 1111001
86 111101000
157 111101001
164 111101010
170 111101011
159 111101100
88 111101101
127 111101110
161 111101111
120 11111000
87 111110010
163 111110011
19 1111101
51 11111100
129 111111010
155 111111011
17 1111111
vinicius�}���T��l^~^~���g�����'��'+ri[�JܚV�_���#?r3�#?r3�#?r3�#?r3�#?r3�#?r3�#?r3�#?u����_���Y~�/�e���u����_���Y~�/�e���u����_���Y~�/�e���u����_���Y~�/�e���24�24�24���������~�h6��k(6���߼���W8�s�x=�/�W:����UΡ�Ľ5��ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�y7�&��߼���~�o�M�ɿy7�&��߼���~�o�M�ɿx����_�K��~�/�%�ī�B��+�B��+�B��+�B��+�D�D�D�D�D�D�D�D�D�D�D�D�D�D�D�D�R5^_��{�_���������VKe�[.��t�ˤ�]%��-�Il�Ke�[.��t�ˤ�]%��-�Il����k���k���k���k��9}���9}���9}���9}���9}���9}���9}���9}�V�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�Jܺ���\��r��9{�D�D�D�D�B��+�B��+�B��+�B�ī�J�ɫ���ɫ���ɫ�J�Ŀy7�&��_�K��~�/�%�ĥn�+u	-�IlJ�ɫ���ɫ�����dk����f��뜚�ɫ�M�l����dlpl����Ւ�:<��}]������\��+~W�ߕ��w��_�����?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��?`��1�A��|�c�$� ��>J��x�� ��>H1�x�@���>H1�A��|�c�$�<k���k���k���k���k���k��8����:<��<������8����8����8����<C��<C�� ��>O��}�?`��?`��?`��?`��?`��?`��?`��?`���/>�/>�/>�/>�/>�/>�/>�.���P���P���P���P��._��._��._��._��._��._��._��._��4�ɥnM+ri[�JܚV�ҷ&�rj�&�rj�&�rj�&�rj�&��_���Y~�/�e���u����_���Y~�/�e���u�di��4��pl�86F�#N���Ӄr�7(�r�7(�r�7(�r�7(�r�7(�r�7(�r�7(�r�7(��ܐ��ܐ��ܐ��ܐ��ܐ��ܐ��ܐ��ܐ��L���L��@�*�P6/?/>?>??P��3������4�ɥnM%�g����܌���܌���܌���܌���܌���܌���܌����e���u����_���Y~�/�e���u����_���Y~�/�e���u����_���Y~�/�e���u����_���Y~�/L�?L�?L�?L�86��k/�M�ɠ��������y7�&��߼�ٔ��*��fR���}s�W:�s�A�9��9��9��9��9��9��9��9��o�M�ɿy7�&��߼���~�o�M�ɿy7�&��߼���~�/�%�Ŀx����_�K��~�/�%�Ŀx����_�K��~�7��7��7��7��7��7��7��7�:��:��:��:��:��:��:��:��݂����h�:��:��k4`ܝ�[�Il�Ke�[.��t�ˤ�]%��-�Il�Ke�[.��t�ˤ�]%��-�J݂V��`����%n�+v	[�JܺV�ҷ.��t�˥n]+r�[�r�/�r�/�r�/�r�/�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�ImD䶢r[Q9-����NKj'%��ډ�9{뜽��^��Q:�Q:�Q:�Q:�Q:�P�u
�P�u
�P�u
�P�q*�&�rj�&�rj�&�rj��q/�M�ɿx����_�K��~�)-�IlJKbU�M\�ߺ��u���3��.��5�l�|#_����Y��:�|#c�dlpl���a����['G��O�˹}���9k���o��[�V�.��+�n�}^}^}^}^}^}^}^|~���~���~���~���~���~���~���~���~���~���~���~������^���^���^���^�>H1�x>׃�A��|����^���^���^���^���^���^���^���^���^���\~���^}^}^|~���~���~���~���c�$� ����^���~���~���~���~���~�������������������������������������������������]������������&��4�ɥnM+ri[�JܚV�ҷ&��4�ɥnM+ri[�JܚV�ҷ&��4�ɥnM+ri[�JܚV���M\���M\���M\���M\�ߺ��Y~�/�e���u����_���Y~�/�e���u����Pl�86F�#N���Ӄdi��4��pnQ�nQ�nQ�nQ�nQ�nQ�nQ�nQ��!���!���!���!���!���!���!���!���!��!�`�@�<��C��8�L��L��L��L�|JV�ҷ&��4���KH��e���������������nQ�nQ�nQ�nQ��~�~�~�~�~�~�~�~�~�~�~�~�~�~�~�~��Ӕzr�NQ��=9G�(����Ӕzr�NQ��=9G�(��,��,���~�pme�Pme�Pme�Pme�Pme�Pme�^�"_�$K��ʾ̥Mf��%\�Ρ�����������������ɿy7�&��߼���~�o�M�ɿy7�&��߼���~�o�M�Ŀx����_�K��~�/�%�Ŀx����_�K��~�/�%�Ŀx����_�K��~�/�%\�Ρ\�Ρ\�Ρ\�Ρ��P�3/L������0���<��\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'+v	[�J݂V��`����%n�%��-�Il�Ke�[.��t�ˤ�]%��-�Il�Ke�[.��t�ˤ�]\�Ρ\�Ρ\�Ρ\�Ρ\�Ρ\�Ρ\�Ρ\�Ρ\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'\�'����������������Ŀx����_�K��~�o�M�ɿy7�&��_���Y~�/�e���y7�&��߼���~�o�%�Ŀx���q7�8��y;�����N�Y��h���>���F�鑪�dj�mf�Y���������686F���f�r�r4���������[�JܺV�ҷ.��	�m�䷶��ݕ�	�yy�yy�yy�yy�yy�yy�yy���q��q��q��q��q��q��q��q��q��q��q��x>׃�x>׃�x>׃�x>׃�A���������ϣ�Ϗ�<j|����^���^���^���\~���~���~���~������\~���~������������~���~���~���~���^���~���^}^}^|~���~���~���~���^}^}^}^}^}^}^}^|���_Q/����_��/������}D�}D�|K�Ĺ|K�Ĺ|K�Ĺ|JV�ҷ&��4�ɥnM+ri[�JܚV�R��������me+k)[YJ��V�R��������me+k)[YJ�ʹɫ���ɫ���ɫ���ɫ���Y~�/�e���u����_��� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܢ� ܣ�L���?M2~�d�4��i���'�N� ��� ��� ��� ��� ��� ��� ��� ���Zx�Oi�*�P6/?/?P��3��3��3��3��3��4�ɥnM%�3�ՙ�i�����������������nQ�nQ�nQ�nQ鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧鑧��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�NQ��_��_��_鑧鑧�Pme�Pme�Pme鑧鑧鑧鑧鑧�ī�BKe�Ρ�Ľ5��5��ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�����������������������������������������������������~�/�%�Ŀx����_�K��~�/�%�Ŀx����_�K��~�/�%�Ŀx����_�K�Y�⑪�:�����W:���j����Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q9-�Il�Ke�[.��t�ˤ�]%��-�Il�Ke�[.��t�ˤ�]%���Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�P�u
�P�u
�P�u
�P�u
�P�u
�P�u
�P�u
�P�u
�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q?�&��&��&��&��&��&��&��&�7'v���݃rs�rs�rs�rs�rs�rs�rs�k(6��k(6��k(6��dd# ���6FA�2���������������������уk4`��6�G�#U���|YIR_�L���K����,���F�鑪�dj�nN��)�Ӕ��Z�r�r5Y-��+q7�yt��NKj'%��ډ�:��9{뜽��^�[��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G���q��q��q��q��q�G��/����_�����~���~���~���~���~���~���~���~���~���~���~���������/���yy�yy�yy�yy�yy�yy�yy�yy�yy�yy�yy�yy����}E����[����������������������������������������������������/������}E����_Q/����O�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|JV�ҷ&��4�ɥnM+ri[�JܚV�R��������me+k)[YJ��KH�-#$����2KH�-#$����3�Y~�/�e���u����_���Y~�/�e���u����_��� ܢ� ܢ� ܢ� ܣ�L���?M2~�d�4��i���'�O�L���?M2~�d�4��i���'�O�$_�/�I����RE�)"�����kH6��kH6��kH6��kH6��kH6��kH6��kH6��kH6��V�*��Zx�OP�5P��3��3��3��w�y;�nM+ri[�JܚKH�-#$���r��r�7(�r�7(�r�7(�r�7(�r�7(�r�7(�r�7(�r�7(����Ӕzr�NQ��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�NQ��=9G�(��/�����H�d��H�e⬼U��F{$d/��/��������w�Y~�ޡ⬡|��R�e쑧쑧쑧쑧쑧쑧쑧쑧⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e���œ��'?N~,��Y9��s�d��Ľ8����^�KӉzq/N%�%띂�<1�~�87P�v��/�n��n��n��n��n��n��n��n��n��n��n��n�\�Ρ\�Ρ\�Ρ\�Ρ�Ŀx����_�K��~�/�%\�Ρ\�Ρ\�Ρ\�Ρ�Ŀx����_�K��~�/�%�Ŀx����_�K��~�/�%�������������������PnNpme�Pme�Pme�Pme�Pme��6FA�2��nQ�nQ�nQ�l�86F�#N���Ӄdi��5�l�|#_���dj��̿�F�⑰�2���K^̥�fR�/L��1�2���K^̥����#a�H�}9Lޜ�oM2צ�j�K�5�2�&��*�&�rj�&�ro�%���������%��ډ�mD䶢r[Q9-����NKj'+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+v��	�݄�n�r�a9[����NV�'+v��	�l��΢�s��%���݄�n�}^}^}^}^}^}^}^}^|~���~���~���~�������R�a9[����NKe��{�^�[����NV�'+v��	�݄�n�r�a>�.����������n&�[��V�o���.���.���.���.����������������������������������4�ɥnM+ri[�JܚV�ҷ&�ՙ�j��frZ�9-Y����KVg%�3��2KH�-#$����2KH�-#$����2KH�-#$����2KH�-#$����_���Y~�/�e���u�di��4��pl�86F�#N���Ӄr�6��i�6��i�6��i�6���L���L���L���L���L���L���L���L��S����O���?e>~�|����)�kH6��i�6��i�6��i�6��i�6��i�6��i�6��i�6��V�*��Zx�OP�5?>?>?>�'G���ɥnM+ri[�Ij�䴌�r��r��r�7(�r�7(�r�7(�r�7(�r�M2~�d�4��i���'�O�L���?2~*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?}2�}2�_)8_)8_)?d��H�d��V^�쑐�R~�e��"�rH��Q�T|�$<��e�d�8_)��w�Y~�d�?d�?d�?d�?d�?d�?d�?d�?d��H�d��H�d��H�d��H�d��H�d��H�d��H�d��H�d�?d�?d�?d�?d�?d�?d�?d�?e⬼U����V^*��Yx�/N~,��Y9��s�d����œ��'?N%�Ľ8����^�KӉzq(^F�����?�O��I��J<����}8����^�KӉzq/N%�Ľ8����^�KӉzq/N%�Ľ8����^�KӉzq/N%�ī�B��+�B��+�B��+�B��?x����_�K��~�/�%�Ŀx����_�K��~�/�%�Ġܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�5��5��5��5��5��5��5��24�24�9G�F��(������~�~�~�~�~�~��Ӕzr�NQ�O�L���?M2~�d�4��r��r����|T˾*e�2G�L��Q�e%��K^̥�fR�/L��1���~�#7�H��3{�н3/L��1�2���K^̥�NS7�H��1�i�`ܤ�s#_+rn_&�rj�&�rj�&��_�K��~�7�mD䶢r[Q9-����NKj'%��ډ�ܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�JܺV�ҷ.��t�˥n]+r�[�J݄�n�r�a9[����NV�'+v��	�݄�n�r[/}s��\�.�l��a9[��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��G��/�J݄�n�r�a9-��Ke��{�E�[����NV�'+v��	�݄�n�r�.���_Q>_Q>_Q9[��V�o����N�G�tywG�tywG�tywG�tyw/��/��/��/��/��/��/��/�����+q7��M�|���+q7��M�&�ՙ�j��frZ�9-Y����KVg%�3�ՙ�j��frZ�9-Y����KVg%�3��2KH�-#$����2KH�-#$���r��r��r��r��r��r��r��r��di��4��pl�86F�#N���Ӄdi��4��pl�86F�#N����d�2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�$=2C�O���?e>~�|����)��S����zc�Lu鎽1צ:��^���zc�Lu鎽1צ:��^���O{)�e=짼C��8�K�ĺ<��ɥnM+ri[�J��KH�-#?u�#N� ܣ�L����S*c�Lx��1�<TǊ��S*c�Lx��1�<T�����S'�O�L���?2~*d�T�����S'�O�L���?2~*d�TǊ��S*c�Lx��1�<TǊ��S*c�Lx��1�=���������|��|��|���3�#<U��F{$d/��rH��Q�֨���hV�N����L��Y{��$�����!|��|��|��|��|��|��|��|���3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#<U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬽8�����ʲLz2I�Fw)�d���Ľ8����^�KӉzq/N%�Ľ8����^�KӉzq/N%�Ľ8����^�KӉzq/N%�ī�B��+�B��+�B��+�B�� ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�y7�&��߼���~�o�M�ɽ24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�24�T����2~*c�L����S'�O�L���?2~*d�T�����S'�O�$_�/�I����T˾*e�2w�$Q�I}�E_d�W�$U�I}�E_e3�H��h�S4{$�~�#�/Z���W�j��\B���d���$s�I�T�*f�3G�H��1���~)"����dk�f|�M���r3�#?u�YA��YA�9�lJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�ImD䶢r[Q9-����NKj'%��ډ���ˤ��u�&��|��NV�ܾ���'��'��'��'��'��'��'��'���]���]���]���]+r�[�JܺKj'%��ډ�8��M�[Q9-����NKj'%��ډ�mD䶢}]���%��\�%+ri[�Jܛ�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|K�Ĺ|JV�ҷ&��4�ɥnM+ri[�Jܚ����r��r��r��r��r��r��r���2KH�-#$����2KH�-#$����2KH�-#$����2KH�-#$���r��r��r��r��r��r��r��r��di��4��pl�86F�#N������/��/��/��/��/��/��/��'�O�$=2C�$=2C�$=2C�$<U����V�*��Zx�Oi�<U����V�*��Zx�Oi�!x��x��x��x��x��x��x��x��1צ:��^���zc�Lu鎽1צ:��^���zc�Lu鎽1צ:��^����8�L��K�ĺ<��ɥnM%�3������ZFIi�Ӄdi��D�x��1�<TǊ��S*c�Lx��1�<TǊ��S*c�Lx���S'�O�L���?2~*d�T�����S'�O�L���?2~*d�TǊ��S*c�Lx��1�<TǊ��S*c�Lx��1�<TǾ�����|/��/��/���F{$g���H�_)?}2��w�Z��Հ���o7��}s�Im��#>u�>�e�*��N�N�N�N�N�N�N�O�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�#=�3�Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*�œ��zq/ef�ef�N%�,��8����^�KӉzq/N%�Ľ8����^�KӉzq/N%�ļY9��s�d����œ��'?N~,��x����_�K��~�/�%�Ġܜ�ܜ�ܜ�ܜ�ܜ�ܜ�ܜ�����~�o�M�ɿy7�&��߼��#O�#O�#O�#O�#O�#O�#O�#O�#OӔzdi�r�L�?NQ鑧��=24�9G�F��(������~���Lx��1�<TǊ��S*c�L���?2~*d�T�����S'�O�Z��]�V��$�>�"��H��(�$�>�|�����O���������}��>��?d���$s�I��G8^�q֮=����X^�q֮!z�ǲH��9�$�~*f�3G����$c�I�RE�6�G���%�d���r3�#?r3�# ��Pme�U�M\���M\���M\���M\��[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[Q9-����NKj'%��ډ�mD䶢|��+r�-����NKj'%���w/�r������������������������ywG�tywG�tywG�tywG�JܺV�ҷ.�ډ�mD䶢u�&��|��NKj'%��ډ�mD䶢r[Q9-�tz�G�tz�/�r��/�JܚV�ܾ%��\�%��\�%��\�%��R�&��4�ɥnM+ri[�JܚV�ҷ&��4�ɥnM+ri[�JܚV���Ru�Ru�Ru�Ru�Ru�Ru�Ru�RrZFIi%�d���ZFIi%�d���ZFIi%�d���ZFIi%�d����Ru�Ru�Ru�Ru�Ru�Ru�Ru�Rpl�86F�#N���Ӄdi��4��~����������������������d�4��d��Hzd��Hzd��Hzd����V�*��Zx�Oi�<U����V�*��Zx�Oi�<U�/�/�/�/�/�/�/�/��:��^���zc�Lu鎽1צ:��^���zc�Lu鎽1צ:��^���ty7G�ty7G�Ii%�d����Ru�Ru�R������5
 6�d��Id��Id��Id��I�e����^�8^�>�v�H~�/|���|���|���|���|���|���|���|���|��֞���Z{�O}i�=��/$;��J�Ӗ��庰*�r��䇾H{䇾H{䇾H{䇾H{�/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB�ǾH{䇾H{䇾H{䇾H{䇲F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�(�e̣ٔ{2�fQ��=�G�(�e̣ٔ{2�fQ��=�G�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F��F��F��F��F��F��F��F��F��F��F��F��F��F��F��F����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��#=�2�N�N�N�N�!|��zb�N�!|��zb�N�!|��zb�N�!|��zcӔx���Hx�����V��!֧֧֧֮�����}}>���W�O��I|T��*}_j_�O����S��)�}��>��8^������t{�=����>�v�O�ܧ��S��)�{��=���?�/$u�䎰����:��GX^H��az��������I�4�>�~^;k���S���g���V������"�d�|#?u����_���Y~�/�e������ɫ���ɫ���ɫ���ɿu����_���Y~�/�e������ɫ���ɫ���ɫ���ɿu���3��g����Y��?�f���n�+u	-�W97�86F�Ӕ���]�ؔ�Ĥ�%%�)-�IlJKbR[�����%n�+u	[�J�BV��P�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�rj�&�rj�&�rj�&�rj�&��_���Y~�/�e���u�rj�&�rj�&�rj�&�rj�&�Wn 94/Z��Ӯrj�&��^������Y~�/�e���u����^�������������������������d�4��i���'�O�L���?M2pnQ�nQ��d�4�����RE��"��H��(�$�>�"��H��(�$�>*e�2�H�֪�����"���w�$_�/�V�*��Zx�Oi�<U���?e>~�|����)��S����O����S��{�O{)�e=짽�����S��z�������n��n��n���?�~+t�V�����[��N�����^C��way�/!݅�;���w���������ɺ<��ɹz�䴌��2��N��N��N�� ܣ�# ܣ��Њ�m���C�$=�C�$=�C�$=�C�$ ���j~�!��j~�!��|���|���|���|����j}������+S�V�ܭO�Z�r��֞���Z{�O}i�=�����䇾��[���t|2U��}i�|���|���|���|���^���^���^���^���^���^���^���^���|���|���|���|���d��H�d��H�d��H�d��H�_)8_)8_)8_)8_)8_)8_)8_)8^���^���^���^���^���^���^���^���d��H�d��H�d��H�d��H�d��H�d��H�d��H�d��H�d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?d�?e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬼U����V^*��Yx�/e⬽�3�#!|��|��|��zb�!zb�!zb�!zb�!zc�$=�C�$=�C�$=�C�$=���Hx���H{+Oei�нjp�jp�jp�j~�}}>���G��ܧ�����j���/���S��)�ax�^�������z~o|wG�;���ܷ\w-����;����������q��8���w����@��P>�����@��P>��z��p��_���L��(�9I��4�ɠ�c�$+���d���W}9G�F~�g�����e������#?u��F~�/܌��_����u����_���Y~�/�e���u�s�W95s�W95s�W95s�W97�?�f���u���3��g����Y�s�W95s�~�3��g������dk�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�Ĥ�%%�)-�IlJKbR[�ؔ�ī���ɫ���ɫ���ɫ���ɿu����_���Y~�/�e���u����_���Y~�/�e���97��k�$Q��U�M\��l�?NR�6F�#N���Ӄdi��4��pl�?NR�NR�NR�NR�NR�NR�NR�NR�M2~�d�4��i���'�O�L���87(�r�7(��'�O�$_�/�I�$�>�"��H��(�$�>�"��H��(�����j���/܎��Gp����j�/O��/�V�*��Zx�Oi�<U���?e>~�|����)��S����O�/�/�/�/�/�/�/�/����Sмvp�vp�v~�u��u��u��U��U��U��U��U��U��U��U�v�����^C��way�/!݅�T}���u�dv���vV�R��������ZFW9I�9Es�~�g��?M2pm1��?yG�Hw#�}�C�$=�C�$=�C�$=�C�$=�C�$=�C�Lx��d��Id��֞���Z{�O}i�=�����S��{�Ow)��=ܧ���r��֞���Z{�O}i�=�����S���z��U�����������������������������������������������������������������������S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r�����ߔ{�~Q��=�G�(����ߔ{�~Q��=�G�(���|����|����|����|����|����|����|����|����|����|����|����|����|����|����|����|��H�d��H�d��H�d��H�d��H�d��H�d��H�d��H�d��H�fQ��=�G�(�e̣ٔ{2�fQ��!zb�=�C�$=�C�$=�����֞���Z{�O}i�=�����֞���Z{�O}i�=�������^����}>�}>�}>�r;W�O��S��q�?8��>�r;k����B��н?7�;���ܷ\w-��u�r�qܷ\w-�;w��������J�ܷBw-�]�tr�ܷAw-�]�tr���!z|$/O����>��B��H^��]���8O}?��H��a�i�k���|�Kdޚd�2B���l���S��S����Ӕzr�NQ��=9G�(��l��dd# ���6FA�2���~�~�~�~�~�~�~�����~�o�M�ɿy7�&���me�Pme�Pme�Pme�^�~�~�pme�_����~�j�&�rj�&�rj�&�rj�&�ri-�IlJKbR[�ؔ�Ĥ�%%�/�M�ɿy7�&��߼���~�o�M�ɿy7�&��߼���~�j�&�rj�&�rj�&�rj�&�ro�e���u����_���Y~�/�e���u����_���Y~�/}>_�$Q��/��U�M���9K�T˰l�86F�#N���Ӄdi��4��~*e�2w�L��]�S.���|T˾)"���H��$_�/�I����RE��d�4��i���'�/�I��������"��H��(�$�>�"��H��(�$�>�|�r;��n��c�R���ֻ��>��_ejﲟ?e>~�|����)��S����O���?e>~�|����)��S������o������x��v�^;|/����o���������u��*�r�G�n��]�[��-�}���u�e���w�!���u}�_|�W�!���u}�_|�W�J��R��V�>*T��������2KH��):�):�(�r�沃r�i� �b���l����jp�jp�jp�jp�jp�jp�jp�j~�}��!�=�C�$<TǲH{���)��=ܧ���r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ���r��S��{�OB�C�Zw)�u󎻔����䇪��V����Zz�OUi�=U��H|��H|��H|��H|��H|��H|��H|��H|䇪�?Uj~���U���S�V��O�Z��H|��H|��H|��H|�r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��s)>�R}̤��I�2��e'��O���s)>�R}̤��I�2��e'��O����F{�g�F{�g�F{�g�F{�g�F{�g�F{�g�F{�g�F{�g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�F{$g�(�e̣ٔ{2�fQ��=�D/LB��/L{䇾H{�r�>�j~���Z{�O}i�=�����֝�{�Ow)��=ܧ���r��Sмu�P�=����r�r;w���K����8�U�ת�j�f��ٽV�~�w>廟r�qܷ\|�]~t��;w�T��y�R���_�T��+�!�@t���J��Ң~t���*'�J��Ң~t���*'������~��}�߾���|w�;��O��|YN~��oek4/O����S����=�t�r�G�Zx��^�8^�86Fzr�NQ��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�L�?L�?L�?L�?L�?L�?L�86��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k/e2ﲙwŔ��#N��y5s�W8����_���Y~�/�e���u�s�W95s�W95s�W95s�W94YA��YA��YA��YA��YA��YA��YA��YA�����_���Y~�/�e���u����_���Y~�/�e���u�#N���Ӄdi��4��pl�86F��)|#O�Y~�/�e���S.�$�>������������������������*e�2w�L��]�S.���|T˾)"���H��$_�/�I����RE��d�4�����RE����ejﲵw�Z�֪�����j�/Z�֪�����j�/Z����#�~v�_;u������k�������0�v�^;|/����o������x��v�^;|/����o���������u�}���w�n��]�ۮ���ax���u�}���w�J�ܥQ�R���:��*�/J�ۥ�zU^�/Ҩ���x^�G�J�����X}�_}+�C��a�Ұ��8^C��x�y���ZFIi\��Q\��d�4��ܛ��{)������Hx�����S��{�Ow)��=ܧ���r���Way!��v�]��/$ :U��=ܧ���r��S��{�Ow)�v8��q�����g�����;>�=ܧ���r��S��{�Ow)�}i�=��r��S����Z{�OUi�=U����V����Zz�O��������������������������������Ui�=U����V����Zz�OUj~���U���S�V��O�Z���?�������������������������������������������������1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)�~Q��=�G�(����ߔ{�fQ��=�G�(�e̣ٔ{2�^���^���^���^���^���^���^���^���^���|����j}���������)��=ܧ���r��S��{�O|㯜u�q��:��_8��{��}�ܷ_ܷ_ܷ_�]�ۨ����+J�۳@v��V�*��J���}|4�T���R��r$!�xd8/���}��p^�!�t�8ޜ�Ӑ�z�$-��r$!�@r$!�@r$!�@r'���F|�џ;tg���F|�џ:TO�;ܧ��S.=�G8^�����c�Ge�u���^�O7r�F�O�O��$?u��Hx���Hx���Hx���Hx���Hx���Hx���Hx���Hx��NQ��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�L�?L�?L�?L�?L�?L�?L�?L�?e2ﲙwŔ��#N��y7�&�q(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6��k(6FA�2��l��dd# ���NQ��=9G�(����Ӕzr�2~*d�T�����S'�O�L���86FA�2��l���*d��E�j�H��$_�/�I�$���E��"�d��H��$_�/�I�$���E��"�d�|/Z�֮�����j�/Z�֮�����j�H��$_֮�����jﾟG�O���������}>_�O�������}>_�O��Iaz�_}>_��܎�����z�_d�F�х��az}^�F�х��az}^�G������j��}�ھ��_|v��;W�n��[����~�_�n��[����~�_�����[����~�_�J��a�Ұ��X}��>�U�}+��k�J��Z�Ұ�$<}��rC�ܐ�w$<}��rC�ܐ��-�;��>�Ϲ-��2KH��(�r��(��'�O�L�����b���]��g���u�:U��=ܧ���r��S��{�Ow)��v��{�����Sм���W{��r��S��{�Ow)��=ܧ�q�����g�����;?�v8����r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ�U����V����Zz�OUi�=U����V����Zz�OUi�=U����V����Zz�OUi�=U����V����Zz�OUi�=U���S�V��O�Z���?Uj~���rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$>rC�$;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ>rC�$>rC�$>rC�$>rC�$;��r��S�c�Lw)��1ܦ!zb�!zb�!zb�!zb�=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$;���+S�����������g�q��:��_8��|㯜u�=V���[��s�nz��U�ܥ>r�t��:U�T�G�J��a�R��d<�7NC�Ӑ���>�	n�-���?=	�[����e��9n'�-��帞��3�-��-�	n��-�w��=�}�z�c޷��e��c��|2ݏ�[���v>n��-��r$!�@r$!�@r$!�@r$!�KU9gz�c��w)�}����?7����L���-P���:>r_}>��v�H~�/ei�=�����V����Z{+O��I��I��I��I2~*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?L�?L�?L�?L�?L�?L�?L�?L�?R�R�R�L�?L�?L�86��k/L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?L�?NQ��=9G�(����Ӕzr�NQ��=9G�(����Ӕzr�2~*d�T�����S'�O�L���?NQ��=9G��?d��H��$_�/��Waz��^�v�]��Waz��^�v�]��Waz��^�v�]��Waz��^�v�]������}��>�}}>���G�O��х�Waz��^�w�O����Gj�#�{�ڽ���wr;���܎��Gp�#�{��>�"�/Z��������|���/֪�$�>��_|v��;W������j��}�ڽ�t�r�/ܷK�-���t�r�/ܷK�-���t�r�/ܷK�-���t�r�/ܷK�-���t�r�/ܷK��X~t�>�תC���w$<}�rC�ܐ��$<}�rC�ܐ����9o7�[���|��9o7�[���w%�}�o�r[�ܖ��i\��Q\��d�t��d�����e>~������+Oei���J������;?�v8��q�����gҮ��C�n���d�u�[���J��Pu�Pu�Pu�Pu�Pu�Pu�Pu�Pu�Pu�Pu�Pu�Pu� 8��Oz��U=ꧠ8��n@q�@q�@q�@q�z��U=ꧽT����Sު{�Oz�OUi�=U����V����Z@t��t��t��t��t��t��t��t��t��:}�>��|O����������H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��H|��Hz�S�V��O�Z���?Uj~���U��)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S�c�Lz�S�V��O�Z���?Uj~���U���OUi�=U����V����Zz�OUi� :|�:|�:|�1��1��6���۞s�nxm���<6���۞s�nxm���>r�r�RT�G�J��r��j��t�9oGB[��Kw	n�o�ޖ��%���n�-��帞��3�-�w��=�}�z�c޷����=�}���_����������-�~��Oз���?B�'�[��|��o��d;�a��<2��C���v��-��(2.V��J��[�>v�>��ek��G�J�Ӯ����{�}���v�=���1�н=�н=�н=�н=�=�����V����Z{+Oei�O�L���?2~*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?2~*d�T�����S'��NQ��=9G��?2~*d��E�*d�T�����S'�O�L���?2~��Ӕzr�NQ��=9G�(��*d�T�����S'�O�L���?2~*d�T�����S'�O�L���?2~��Ӕzr�NQ��=9G�(��*d�T�����S'�O�L���?2~�"�d��H��$_�/�I�$���E�*d��E��"�^�v�]�I����S'֮�����j�/Z�֮�����j�/Z�֮�����j�/Z�֮�����j�/Z�܎��Gn�#�{�۽����v�r;w��֧������܎��Gn�#�~v�~�wr;���܎��Gp�#�{��=��}>_�O��Gp��־v�]��}>_�O��Gp�#�{��=���wr;���܎��Gp�#�{��=���wr;���܎��Ұ��X~t�?:V�+Ε��J��a�Ұ��X~t�?:VT�k�!ڀ�p���!��Hx��>䇏�!��Hx��>䇏�o����[�z��=V��~�U�G�ߣ�-��K}{��^�ֹ�+����+���L��Hx�Oi�o�ۮ�-��+OM1�)!�����;?�v8��q�����g���n��Lxd:2�>W��xd:>�c�n���8���8���8���8���8���8���8���8���8���8���8���8�J��܀�U=ꧠ8��nt�S��:��:��:��:�Sު{�Oz��U=ꧽT����V����Zz�OUi�=U���������������������������t��t��:|�:}�>~���U���?Ui�O�Zz�S�V����Zz�OUi�=U����V����Zz�OUi�=U����V�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!�9!����U���S�V��O�Z���?Uj}�c�Lw)��1ܦ;��r��S�c�Lw)��1ܦ;��r��S���U���S�V��O�Z���?Uj~���Zz�OUi�=U����V����Z@t��t��t��c��c��c��m���<6���۞s�nxm���<6���۞s�nz�:>����V���9�!���y�2n��qЖ�:�B��-��K�r�z[��[�<6�΄�IӮ����=:폮�_Њ�z��
���_Ю��k���VO-Ed޸���o��k�~��Mз���7B�'�[��|��!�xd;�a��<2��C���výo��ң=Q�/�w�!�xm��9n�-���/��������H��n��K���������/Z�/OB��/OB��/O{+Oei�=�����S����ZB�Ǌ����S�R~*b�O�L{��$����H{��$����H��L���?2~*d�T�����S'�O�YA�2�����L��H��]��W|T�����S'�O�L���?2~*d�9G�(����Ӕzr�NQ��<T����_)?1�'�!|��T�/�������S�R~*b�O�Lzr�NQ��=9G�(����Ӕx���S'�O�L���?2~*d�T��$��H{$��H{$��H{$��HB���������������$������}}>���G�O���������}��0�j�/Z�֮�����j�/Z�֮������^�v�r;W��܎��Gj�#�{�ھ�}}>���G��܎��Gj�����t���k�n��Z�ۭ|�־v�_;u������k�n��c��<����J��Z�ۭw#�{��=���wr;���܎��Gp��־v�_;u������k�n��Z�ۭ|�ֽ��?;u�}+��k�J��Z�Ұ��ֽ��?;u��k�J����ro����-���y�r�o����-���y�r�o����o����[�z��=V��~�U�G�[�ܖ��%���o�r[����!�<U���?e>~�|����;?|v~��������}��q��:��_8��|㯜u�q��:��_8��|㯜u�qת��S�u�^s�nt�S�ҧ�<6���۞s�nxm���<6���۞s�nxm���<6���۞s�nxm���Pu�Pu�Pu�Pu�Pu�Pu�Pu�Puӎ�q�N:��]8�t㮜uӎ�q�N:��]8�t㮜uӎ�q�N�>�uӧϧt����]:|�q�N�>�uӧϧt����Pu�Pu�Pu�Pu�_:��Z|�O�iܒ�!ܒ�c�Zz�OUi�=U����V���ߔ@t��t��)�����o�ۮ��Oi�<5����֞��ZxkN�>}:|�t�������ӧϧO�N�>�>}:|�t�������ӧϧO�N�?i�<5����֞��ZxkH�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�?i�<5����֞��ZxkN�v��v��v��v��v��v��v��v��*}�S�JxiH܀��:�S�8��|�U��_Ү�t��:U����!���z:�}
�^�w�z���]�-T�e��O�ޮ��m�=	n��-�t%�N�V����Wk�qY?z+'�T垸���S�z�n�NM�ɺ97�+gЩɽq[>�VϽS����;�\�O���T�;�<�O�S���l�q[>�vEз���?N[���u�9��!��)Q�	�J��Ҡ`;wX�q���Gq����q�?8���_�O��S���X{�۾�}}>��v���G�����S��{�Ow)��=܎�T�r���}i����$=���H{�O���֟9!�>rC�Z|䇾HB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/LB��/$;��/$;��/$;��/$>rC�Z|䇾���}i����!y!�����^���^��V�ܭO�$]�I{�E��w�$]�V��=�����֞���Z{�O}iܧ���r��S��{�Ow)��=֧�*c�$=��=��_}>�/Z��������U{��~�>_������p�#�{��=���wr;���܎��Gp�#�{��=���wr;���܎��Gp������}�Vn�+7r���!���z>r�T���-���z>r��+7r���n��c�۱����v�;v?���ݏ�n��c��=����@r�C��z 9D!��K|������]�����8^;k���㶽��^�v8^C���w-�=R�8�q�� ;}�o��������@v���q�� ;}�o��������@v���q�p0��p0���mi�<U���?e>~�z�����;?|v~��������_8��|㯜u�q��:��_8��|㯜u�q��:��_8��nxm���<6���۞s�nxm���<6���۞s�nxm���<6���۞s�nxm���<6���۞r��8���8���8���8���8���8���8���8�t㮜uӎ�q�N:��]8�t㮜uӎ�q�N:��]8�t㮜uӎ�q�N:��]8�t㮜uӎ�q�N:��]8���8���8���8���8��Oz��U=ꧾu�δ�I��V����Zz�OUi�=U����S>~��9!�;uޝ�華�֞��ZxkOi�<5������ӧϧO�N�>�>}:|�t�������ӧϧO�N�>�>}:|�t�����֞��ZxkOi�<5���������������������������������������ӧϧO�N�>�>}:|�t�����[����{���u����z�w�n�ޥO�Jw�N���ҞS�J@q�z��U�� :T�:U��w�!��R���9�B[��Kw��w�z�	�������V��]���l;����ýo����:qY?N+'��d�
���S�t*rn�FEިȺ97B�&�El�[>�Vϡ��El�[>�O�S����zu<�W���T�;�<O�S����=q[>�vYз���?N[��Kv=97�-��$8.�+�N�	��Ҡ`;w8�������[�|�`8�;��J�܎�������{�ۿ;u�>�}iܧ���r��Sި��z��Tu�9!�9!�9!�9!�9!�9!�9!�9!��!��!��!��!��!��!��!��!��1��1��1��1��1��1��1��1ܦ;��r��S�c�Lw)��1�=U����V����Zz�OUi�=�����֞���Z{䇾Hw+S�V�ܒ.�$���"�rH�ܒ.�+S�֞���Z{�O}i�=�����S��{�Ow)��=ܧ���r��ۨ��������������V��_��������)���|��;�������p����v�;v?���ݏ�n��c�۱�#����]���v�r;k��܎��Gm{�������Vn�+7�C���|�=�o�/��mB��P�v�/��mB��P�vת���J��f�R�z�Y�T�ުVoU+4!��=����@r�C��z>r��qܖ���=�Gr[��������?�v������o��Wz�qX+������k�|5޾�_w�����]�����z�v���q�� ;}�o��������@r�-��r�-���Oi�=���)�e=�g�g�������۟8��|㯜u�=T����R��S�Jz�OU)�=T����R��S�Jz�OU)޷�޷�޷�Ж�Ӑ�S�J@v熔�ҞS�JxiO)�<4����ҞS�JxiO)�<4����ҞS�JxiO)�<4����ҞS�JxiO)�<4����ҞS�JxiO)�<4�N:��]8�t㮜uӎ�q�B��[�s�nt-΅�з:�N:��]8�t㮜uӎ�q�N:��]8�t㮜uӎ�q�@q�@q�@q�@q׆��ېu�PuꧽT����V����Zz�OUi�=U��������N�w�$>rC�n�ӷ]�V���ZxkOi�<5����֝:|�t�������ӧϧO�N�>�>}:|�t�������ӧϧO�N�>�>~��ZxkOi�<5����֐u�Pu�Pu�Pu�Pu�Pu�Pu�Pu�]8�t㮜uӎ�q�N:��]�T�ԩ��S�R�ޥO�J�z�>�*}9Ӑ�9Ӑ�9Ӑ�:T�t��t��t��d:>�-Հ庰�/�v��}	n�o�з��[�=u߼�g�����jv<�+_����1Y?z+'�Wk�97B�&�Td]ꌋ�Q�z�6~���������8>������ʽu9W��*���]
�B��Щ��*y�
���Q�z�r�]NU��ʽuj�����z�}�싽]�t-�~��ýo��Kt�9n'�!�t$?�:T'NC�Ү :U�n�۳@t�~�u�U�ת�k�n�ܧ����}��?;t���G�O��$;��r��S��{�Oz��TuꎽU����V����Zz�OUi�=U����V����Zz�OUi�=�����֞���Z{�O}i�=�����֞���Z{�O}i�=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�����֞���Z{�O}i�;��r��S��{�Ow)��=ܧ������֞���Z{�O}i�;���+S�V�ܭO�Z�r�>�w�Z�r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ�����W�n��Gj�����k�-��;^�V�>_�O��S��q�?:}�Tw�;����c�۱����v�;v?���ݏ�n��c�۱����v�;v?���ݏ�n�ܥf�R�w)Y�r�����-��K|�R�8^;j���۱�������9G�[�����Y�T�ުVoU+7����J��f�R�xe�~o��[����e�~o��[����m�}U�>��Uw���ܖ���;�|�q���W|�q_�W����xjp��'����]�����z�k�|5޾�_w�����]�����z�k�|5޾�_w�����o��������Oi���O����㳅㳅���g���n{�Ϝu�q��:�R��S�Jz�OU)�=T����R��S�Jz�OU)�=T�����ux1Z>��������?)ې�Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9�<4����ҞS�JxiO)�<4����ҞS�JxiO)ӎ�q�N:��]8�t㮜uз:�B��[�s�nt-΅�ӎ�q�N:��]8�t㮜uӎ�q�N:��]8�t㮜u�Pu�Pu�Pu�PuӥO�J�N�>�*~s�n@q�@t��t��t��t��t��t��t��t��t��)Tz�>���Zt��zv뾪ӧO�N�>�>}:|�t�������ӧϧO�N�>�>}:|�t�������ӧϧO�N�>�>}:|�t�������ӧϧO�N�>�>}:|�t�������ӧ���8���8���8���8���8���8���8���8�nt-΅�з:�B��[�s�J�z�>�*}�T�ԩ��S�R�ޥO�-ϡ-ϡ-ϡ-ϡ-ϡ-Ͻ-��Kwzr�ޜ�w�o��[��6�~���N�k�o�޷���`{�����'+-T�e��l�S���6�F�Z��媜�Z��%���Q�pj2o]��A����84<Z�`�T<�j��-P�%�D�CȖ�y�>Z���T�]?�A���u}t_]W�C�����|�Aϖ�y�"Q�ʥ���Q����=q[?\VM����u�]výo���t��n'�-��$?�T�C�Ӑ���>~V����!��X�:V?�wr;W���a�R����{���������g�8���8���:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|�:|���r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ��C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�C�$=�����֞���Z{�O}i�;��r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ�t��t��t��t��t��t��u�?:}�:}�8��q�����g�����;?�v8��q�����g����Ο����n��Gj�����k�-��;^�V�w�;����Z�Gq����;vhݛ�J��f�R�z�Y�T�ުVoU+7����J��f�R�z�Y�T�ުVoU+7����!���z>r�T���-��K|�;}�o���z=R�8�q����`{���'��	���e�~o��[����e�~o��[����e�~o��[����e�~o��[���{�;�+��Q�Ө����}��mj��������?;|�������>�V����`zqX�V����`zqXw�����]�����z�k�|5޾�_�φ���o����S��{�O{)�^;8^;?|v}�u��S�Jw)N�)�=T����R��S�Jz�OU)�=T����R��S�Jz�OU)�=T����R��N��S������n�%���7����Μ���n����n����n����n����n����n����n����n����n����n����n����o)�<4����ҞS�JxiO)�<4����ҞS�JxiN��з:�B��[�s�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nt-���<6���۞s�nxm΄�BC��!�ӥO�J�N�?�� 8���8���8���8���t����{���:�㮝*}:T�T�N:��]8�t㮜uӎ�q�B��[�s�nt-΅�з:�B��[�s�nt-΅�з:�N:��]8�t㮜uӎ�q׆��۞s�nxm���<6���۞s�nxm���<6�z��R��S�Jw�N�)ޥ;ԧ�C��C��C��C��C��C��C��C�B[�B[�z�z���G�o�ޮ��Wp���{��>��?]wB����ފ��Ey��~}qXNV
Z���U8�F�-Ple����S��5g�&��2)j�g(�p%�A���y�Gٟ��g�m���{JZ�iKQ�)j=�-G�e����Ֆ�ڲ�{VZ�vKV��j����vKV��j��-[;%�gd�Ֆ�ڱ�f��CҔhzR�?�A�ph2�]GZ���U9d�S�pb�]v��]��Wcz�΅v'�-��[��-�zv������-���|�r?���J����[�@t�~o��������[��[��[��[��[�s�n@t��t��t��t��t��t��t��t��t��t��t��t��t��t��t��t�����g�����;?�v8��q�����g�����;?�v8��q��)��=ܧ���r��S��{�Ow)��=ܧ���r��S��{�Ow)��=ܧ���r��S��{�O|���g�����;?�v8��q��㯜u�q��;?�v8��q����������}Q۾���Tv�;w������������������܎��Gn�#�{�۽����v�r;w���K�#�}��=��_U��J��Z��p��}V�^��?Twn�۳@v��V�C��z 9D!��=����@r����-���|�2�?���-���|�2�?T���-��K|�R�8�q��<5޾�_T���-���8�B��Q���phzv�����o����:v�����o����:v�����o����:v�����o����������`8��N�Q�Р�w�q0W������}U�>��UwϪ���S�������j~|5?>��Oφ�����qX+�``8����0V���밐v��{)�e=짡x��x����������r��R��S�Jz�OU)�=T�!�9�hC@r�����4!�9�hC@r�����7+G�]����[��Ks��n���ҝ9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�s�nt-΅�з:�B��[��T�ԩ��S�R�ޥO�J�z�>�*}s�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nxm���<6���۝	���BC��J�N�>�*~s�nxm���<6���۞s�nt$;�5ھ�}��]	��*~�{�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nt-΅�з:�B��[�s�nxm���<6���۞s�nxm���<6���۞S�Jw�N�)ޥ;ԧz��R��S�!��!��!��!��!��!��!��!ϡ-Ͻo��o��]���Ֆ������O����-T�KQ[�]N�Q�����jp2�F
Z��KU8�F����4;	F�_�����Q��%��Q���(x1d�#l�G"��{JZ�iKQ�)F)�(�5c�x�^9 �@;#����9 �@;#�M��Sr9ܖ�۲�{vQ�n�1��F=�(Ƿe��׈ǵ�1�x�V9lՔm���#�A�ph2�j�g(�dҍFM-T����]���l=qZO]�'�o��[�;�����w�z�׽o�Ю���z :V?���-��[��d<ުV���W�J����d:>�B�G�!����������������������������������_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�����;?�v8��q�����g�����;?�v8��q�����g�����;?�v8��q�����g�����;?�v8��q�����g�=V���[��u��u��u��u�*�J�ۨ�v�0��n�ۨ�v�=����v�r;w��܎��Gn�#�{�ۿ;u�����G�n��Q�ۨ���~v�?;t�r;W�O�܎��[�@t�~�u��w��k�n�۳@v��V�+G�����xe�~o��[����e�~o��[������;}�N�qӷ�t��;}�N�qӷ�z��p����@v��w�����]����R�|�=9G�[��� ;}ǆ���]�Ю��Wz�+�z޽
�^�w�B�ס]�Ю��Wz�+�z޽
�^�w�B���]��I}طy*����;|/J�ܖ��(0R�R��l���#;�8��'�C��P`�.��Q�Ө�����?�u�:���G�N���S�������j~|5?>��Oφ�	����~�b�|1_��{�OB��/n{���)ܥ;���C��[@r�����4-�9m�hC@r�����4!�9�hC@r�����4!�9Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ж�Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9Ӑ�9ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)����ޥ;ԧz��[�s�nt-΅�з:�B��[�s�npe��Ȭ��]�ޥO�nz�;�ԩ�iз:�B��[�s�nt-��*}�T�ԩ��S�R�ޥO�J�z�>�*}�T�ԩ��S�R�ޥO�J�z�>��з:�B��[�s�nt-��)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�O\�?\���o\���o\���o\���o\���o\���o\���o\�>�����w�o������mpjx媞�j��Q��j}x5���Q�-T|�5IF�	(�bx4�j�c-Ple�r�'��%���E-PdR�E(�p#�<Fٟ�iDb�����׎@;#����#݈÷b0��$:��qD`QF��qDb�(�R��\����c�R�{�Q�qJ1M�F)�(�7#�M��Sr9 �b���f��CҔhzR�"Q��J4	j�g��ɽu9g��'��k�5;�v7���E~�"����'z���]�ޮ���a:޽;}�N�q����z�~o!ڀ�9~��/Ӑ��r�N[�Ӗ��庰*�J�Ү�t��*�J�Ү�t��*�J�Ү�t��*�J�Ү�t���s�nz��U��=V���[��s�nz��U��=V���[��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u�8��q�����g�����;?�v~�s�nz��U��_�_�_�_ۨ�v�0��n�ۨ�v�0��n��K����;t���/�K����;t���/�K����;t���/�K����;t���/�c�ۭw#�~v�P���-��=;v?U+7����n�Ү :U�J���}|2_���!��H}}R_T���!��H}}R_�φ���o�������m�|6�>�[���[�����m�zu��:���w��C�����>����C�����>���N���]�Ӯ������u��:���w�N���]�Ӯ������u��:���w���Z�J#��b�}����W_�������Rpm��e'��ޠ�w�1�
�OB�Ө���~��?zu�:�ޝG�N���Q�Ө���~��?zu�:�ޝG�N���Q�ө�t�p]:�N�짡x��{r�;��r��R��S�-�r������4!�9m�hC@r�����4!�9�hC@r�����4!�9�o)�:r�!�����������������������������������������������������������r�!�r�!�r�!�r�!�r�!�r�!�r�!�r�!�ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ=r�ԧz��R�s�nt-΅�з:�B��[�s�nt-΅�-[��jxc�Y~�*}s�!�ޥO�Ot-΅�з:�B��[�s�nw�S�R�ޥO�J�z�>�*}�T�ԩ��S�R�ޥO�J�z�>�*}�T�ԩ�-΅�з:�B��[�s�nw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�!�r��-�r��-�r��-�r��-�6��m������σo��>�||�������]���W�S�-TsJ5r�G��S�����>e���F�	(�a%��Q���c%���A��hv��#l�J6��l�KT�A�J4	F=*�G��1M[$^9 �@;#�Ȍ;v#ݲC�,���$:�d�\��땒r�C�VHݒ�d�m� q�r)r�E.Qȥ�9�G"�(�R��qG QF��nJ1Mx�{^9lՔhzR�JQ�ʥ�A���6|���S�KU9g+_޷������gz�����a=qXN�w��Q���a:�=
�^W�+��]��[���;~n����o�޷��[�w�����0*�J�Ү�t��*�J�Ү�t��*�J�Ү�t��*�J�Ү�t���u��s�nz��U��=V���[��s�nz��U��=V���[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[��[���g�����;?�v8��q����[��[��s�nz������������iU|4��U_*���W�J��U�Ҫ����;t���/�K����;t���/�K��X}T�>�VU+����J��a�R��e����J��y�v�}
��N�q����Y�T��*��\@t�����!���}}R_T���!��H}}R_T���!��H}|6�>��φ���o�������m�`9n��|6�>��w�N���]�Ӯ��Ea:XN�V�]�Ӯ�����m�`9n�]�Ӯ������u��:���w�N���]�Ӯ������u��:���w�N�����u�밝�g������1�
�Oz�ޠ�t*1=:��+����a :�'N�Ө���~��?zu�:�ޝG�N���Q�Ө���~��?zu�:�ޝG�N���S����u8.�N�nw)N�)ܥ>r��-�9���hC@r���9mӖ�9mӖ�{�oxm��᷼6������{�oxm��᷼6������{�ot-з��B��[�{�ot-з��B��[�{���S�ޮ��!�:S�!�rۡot-з��B��[�{�oz��������oU�ҞӖ�9mӖ�9mӖ�9mӖ�9mӎ�q�B��R�n��V�
�jS���R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz���w�e��2��n��[��-������s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��o\���o\���o\���o\���o\���o\���o\���o\���R�Nqʍ�Nr�Uޖ�	���5�����j*���F�9F+w�o��o�ޮ���e�5<r�G7��Z���4��r��9A��h11�dr����T��A���ryF�"�G����{Q�J���9҈�5b1�x��#݈�8���Fr�C��W>JϒS�ߒ~;d���N��)��e;��s��}��϶S���w>�?�#���c����?�Q�m�`qݒ�d���!�qu�# �E7#�M�F)��iJ6��Fٟ-[0x4<�Z�ȥ���Q���6���I����p]�ބW�+���pb�^��'�+	ފ����=�^���B�ϡo�ӷ��Ky���n����-��Kxz�����-���r�9_�J��U�Ҫ�iU|4��U_*���W�J����庾��C����t��*�J��_Ү�t��*�J�Ү�t��*�J��݀��`;u�G�J��U�Ҫ��9*���W�J��U�Ҫ�iU|4��U_�����G�n��Q�ۨ���~v�?;u�����V���2������T��:U��G�!���t|2*���W�J��U�Ҫ�iU|6�>v��݇�n��a�[�z�ֽV�^�u�U�ת�k�n��Z��X�:V8���c��X�:V8���c��=����xe�~o�N�qӖ�zr��C�������Ӑ��%��	o�B[�������m��6���������o��~|6�����N�	Ӯ�t밝�ޝv�]���a:u�N�v�]���a:u�N�W�B+���Њ��E~�"�z_��ޝv�]���a:u�N�v�]���a:u�N�N�S��T��8.�N�S��T��8.�N7�S��T�z8ޅN7�S��T�z8ޅN7�S��T�z8ޅN7�S��T�z��F'�Q��Tbz��F'�Q��Tbz��F'�Q��Tbz��F'�Q��Tbz��3�A��Pc;���)ܥ;��r���o����s��s��4-�9m�n����n����o�᷼6������{�oxm��᷼6������{�oxmз��B��[�{�ot-з��B��[�{�ot-���[�������-��-Th����WgޮϽ]�z�>�v}���������Wgз��B��[�9mӖ�9mӖ�9mӖ�9mӖ�9mӖ��S�Jw�N�)���k�b59{%Gz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧz��R��S�Jw�N�)ޥ;ԧ[��-������w�e��2��n��C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�C�[z差[z差[z差[z差[pm������σo��>�||�6����u(����(��-E^�{�-�5�����j*���F�9F�>N﮻w�o�ޮ���e媎iF��Z���U1�$r��9A��Pbc���69A��hv���A���ryF�,�G���8�{Q�`�"����F)��k� �v�r�C�VH~ݒ�B��P�|�������+Կ%z����$�v�?�O����$�~I?�/��%϶�s�\�b0���~9�C�,��J?~�߲C��0땒r��8��M��Sr9lՎG����)Fٟ-P�84<	F��-Pd\���Q��U9?�c��z�q��gz�-T�x1X.V����~�Ⱎ��'z+޷��Wn:�}?]��z[�ޖ�w����o7z�k�-��Kxz���/Ӑ��r�NC���r�9_�!���9~��/Ӑ��r�NC���uzr�_�G�!р�W`:U��v�]��W`:U��v�]��W`:U��F�Q���`8쿆�W�n�Ӑ��t�]9_�J�Ӑ��t�]9_�J�Ӑ��t�]9_�J��U�R���U}T���U_U*���W�J��U�R���U}T���U_U*���W�J����iU|4��U_*���W�J�Ӑ��t�]:U��*�N�k�J�ӥZ�ұ�t�p+J�ұ�t�p+J�ұ�t�p+J�ұ�t�p+J�ұ�r�C����e�};}�N�qӖ�zr�N[���p=9n�-��%��	o�z�	޷�xm��6���������o�������m��6����v�]���a:_��ބW�B+���Њ��E~�"�z_��ބW�B+���Њ��E~�"�z_��ޝv�]���a:u�N�v�]���a:u�N�N�S��T��8.�N�S��T��8.�N7�S��T�z8ޅN7�S��T�z8��F��Q��Ti;�N�F��Q��Ti;�N�F'�Q��Tbz��F'�Q��Tbz��3�A��Pc;���3�A��Pc;���3�A��Pc;����Hn���hC@r�oxm��᷺�B��[�{�ot-��᷼6������{�oxm��᷼6������{�oxmз��B��[�{�ot-з��B��[�{�ot-�U������q[�q[�5;����=k�]�z�>�v}���������WgޮσS�з�:S�-�5;����w�ot-з��B��[�{�ope��2���~�~�rվ�]�����s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��n���n���n���n�������������n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n����6�����{�oKUԵ]KUԵ]KUԵ]KUԵ]pk�j*�js�To�js�js��^�zZ����Z����Q��Q��9Q�Z����h���}q[\�?]OD�A���02��r��#C��P�#�؍�#A���l#�9<r�'�m�.�E-G������E2#�L��SV9 ׎@;"0+$:�d�\�P�J;��߲|p�>8hU.�N�)ԡRL!$��L!$��MJ$ԡ�MJ$ԡ�MJ$ԡ����R�D~?"?����϶�s�\�l�6O�?~�߲C�"0��R��qG"���S^Q�k�Q�)Fٟ-[0e�f�g�Ƚt97�,��l;�;�F��S��T�}u8�]N7�S���bx1X.O�+	���E`z޽�^�v�o�з��[��+�=v��~�����-��Ky�>����!��Ky���n����-��Ky���n����o�Ж��%�=9_�!���9*���W�J��U�Ҫ�iU|4��U_*���W�J��a�۰�mֺt�]:V>�*�BC�А���X�t�]:V>�*�N���J�ӥc�ҭ@r�C��v�9�!ڀ�;P�j��xe�p�k�J��K�����VC�����V�r�N�k�J�ӥZ�ҭt�V�t�]:U��+N���J�ӥc�ұ��X�v���7����J��f�R�z�Y�T�ުVhC��z 9D!��=����@r����!���}zr�N[��[��-�z�=9�NC�Ж��%��	o�z�	ޖ���N���;|o����P�
��@v�/T����@v�(����k�>�O��Ю��+�=
�OB�Ю��+�=
�OB�ފ�w����gz+ފ�w����gz+���k�>�O�����k�>�O��Щ��*q�
�oB�Щ��*q�
�oB�ި�w�4��'z�Iި�w�4��'z�Iި�w�4��'z�Iި�w�4��'z�IӨ�t�4�:�'N�IӨ�t�4�:�'N�IӨ�t�4�:�'N�IӨ�t�4�:�'N�IӨ�t�4�:�'N�Iܐ����9m�o�?�᷼6����[�{�ot-з�u�����gӮϧ]�N�>�v}:��u�����gӮϧ]�N�>�v}:��������WgޮϽ]�z�>�v}���������WgޮϽ]�z�>�v}���r۽]��w�S��������4�f�v}���������WgޮϽ]�z�9j�G�-�V�N[G(r�(�9F�W�ot-з��B��[�{�oG"�e���C��C��C�[��-�������������������������������������������������������������������������������������������������m���m���m���m���վrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվrվr�u-WR�u-WR�u-WR�u-WR�u-WR�u-WR�u-WR�u-WR�U-ER�Nr�Nr�Nr�Nr�Nr�Nr�U(��(��(��������(�j�QY\V_�S�-TsKT�F��9C��P~�-��KdlF�I��Y(u�J��l�Dm���z�9��b��S9�D`Hv����vDa۶Huʅ۔�|��ϒI���w>K��R����M.+���.����{�Xok��a��\�K���q��.?ߥ������K��t���K�P��
!d�B�:�*S�B�8?�
��$�v�w>?~�߲C�,��H��# �E7%��F=��iJ6��F=*���<��C���rnY��z�6�$�A���i85NF�Z���U8�j������a=u?>������������z�q���pk��v�~�~�]��z[�ޖ�w��޻?]�G����o������z���v��o7z�k�o�Ж��%�=9_�!���9~��/Ӑ��r�NC���r�9_�!���V�t�}:V>�+BC�А�w���oGz[�ޖ�w���oGz[�ޖ�w���oGz[���xe�~7�[���xe�~7�[�Ӗ�xe�~�u���_���a��y�v��	BC�А��$<}	BC�А�t$<��oGz[�ޖ�w����zC�ސ���>}9��[����e�~o��[����e�~o��[����e�~o��[����e�}9n�-������B��o�ޮ��W�%��	o�B[�޷�w����]�'�]���b|5؟v'�]���b|5؟v'�]����P��]���b|5؞�V3����c;�X��V3���Ec;�X��V3���Ec;�X��V3���Ec;�X��V3���Ec:qXΜV3����c:qXΜV3����c;�N�F��Q��Ti;�N�F��Q��Ti;�N�F��Q��Ti;�N�F��Q��Ti=t]��A���l}t]��A���lzuN�F��Q���i:uN�F��Q���i:�ǡA��Plz�ǡA��Plz�ǡA��Pl~r��-�r��oxm��Ӯϧ]�B��[�{�ot+��uЮ��N�>�v}:��u�����gӮϧ]�N�>�v}:��u�����gӮϧ]�z�>�v}���������WgޮϽ]�z�>�v}���������WgޮϽ]��vZ�юP�媍\V��v~����F��+�+�+�+�+�+�+�+|�A�з�V�N[G(r�(�8�_�]�B��[�{�ot-з��r�FQ�ݖ���m���o\���n�~�m�޹m�޹m�޹m�޹m�޹m�޹m�޹m�޹m�޹m�޹m�޹m��m���m���m���m���m���m���m���m���m���6�����{�opm�j����j����j����j���������rގ[��z9oG-������rގ[��z9oG-������rގ[��z9oG-������rގ[��z9oG-�j����j����j����j����F*�b�F*�b�F*�b�F*�b�F+vQ�ݔb�e��F+v9S��ղPe���F+v9S��юT��j5b5����S�-TsKU��9F��9l��}��଑�K%���C��[$�+d��C�Jv�;%��#��E%QȤ�# ȲC��P�X�;��ݡ\��?��
��)�o�?�O�l�R�J�(T��J���K�w���g��x�x��X�xՈ��X�xՈ��N�x�跍N�x�跍N�x����)񭲿�+�N�?$�c�N�)��L!$���J)ԡT*�m��S��С��(w%�r�C�Qv�r��k�1MYF�(ǥR�{Z�`pm�)F�"��r~��A��h5��Z��KTj�c���J5�F��������U?���WϮ�����>���+��]��Wn;������B[��[���>��_]v������}u�\W��ߣ�o����Ky���n����!��Hx���n����-��Ky���n����-��Ky�n�+GzC�ސ���>~�n��-�z廏\�q��=r�Ǯ[���w�n��-�z廎��qз��Kw>��qз��Kw>��qӖ�xiZ<2o+G�C�Ӑ��-���ގ����-��Kz;�ގ����!��H|�r�Ǯ[���w�n��!���8\�Ж�z�N[���p=9n�-�����Ӗ�z�=����B��o�з��[��-�`9n�o�������밝:�'N�	Њ���a:u�N���]��Wbz؞�V3����b|5؟v'�]���b|5؟v'�]���b|5؟v'����c:8ޅN7�S����}u8�]N7�S����}u8�]N7�S����}u8�]N7�S����}u8�]N7�S��Ti;�N�F��Q��Ti;�N�F��Q���l}t]��A���l}t]��A���l=u]F��Q���l=u]F��Q���k�4���A���k�4���A��Plz�ǡA��Plz�ǡA��P�;�;�ýC��P�;�;�ýC��Plz�ǡA���o���[ޫ{�ot���gӮϽ]w���uޮ��Wz*�E]諧t���gӮϧ]�N�>�v}:��u�����gӮϧ]�N�>�v}:��������WgޮϽ]�z�>�v}���������WgޮϽ]�z�>�v}��媍F�V9C��h5}q[��z�?\V�\V�\V�\V�\V�\V�\V�\V�\V�j�G�]�N[t-�j�F9C���4{������WgޮϽ]�z�>�v}������*te��j��[z差[pm������σo��>�||�6��m������σo��>�||�6��m������σo��>�||�6��m����-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-[�-WR�u-WR�u-WR�u-WR�u-WR�u-WR�u-WR�u-WR�u����rގ[��z9oG-������rގ[��z9oG-������rގ[��z9oG-������rގ[��z9oG-��-WR�u-WR�u-WR�u-WR�u(�R�U(�R�U(�R�U(�R�U�єb�e��F+vQ�݈�jШxe;e��N�r�F9S��Ո�j�(2�J�r��9Q�(�tG(|�4>��g��z�l��G�(Q�
zl��q�4�l��c�L{���@2"0�$;>�ҡC�e;��
�B��I5-�&��$Ըex?o~
���P�.�����7����<h�[���u�@{�������}1M衊oEH=1 �Pă�CEH2�{��o~��>�t3�C>�wyX��#����������^�@�`�	N�)��$���'�S���p��?n�۲C�Qv�r��k�`�ȦDr)*�c�1����l�J6�d�l�G(rx�O(�k�|�C���61�lr�-T�e���Q���e���j���������|�b�x1_>���������{�����������>��������<���σ]�������z��=v��o7�ߣ�o������z��=v��~�]��zC���=r�Ǯ[�����m�x6��^���׃o��������m�x6��_]v�]���`}u�]v�]���`}u���q޷���`x1_<��]v�o�Ж�=v�~�?]������-�z廏\�q��86��^��-���~x2ߞ��o�޷��[��-�z�=����B��o�ޮ��W�����������w�z���]���������u���ބW�B+���Њ��E~�+�=
�Oz+ފ�w�����oN+ӊ�tⱝ8�gN+ӊ�tⱝ8�gN+ӊ�tⱝ
�oB�Щ���4��'������q���o������q���o�I���pj4��'�I���pj4��'��c����6>����c����6>����c����6>����c����6>���_����h5��_����h5�|�C��T9<�C��T9<�C��T9<�C��T9?z�aޡ�w�v��z�aޡ�w�v����_�W����e��_�W����eB�cР��(6=
��[|巆����:��u��⮜Uޮ���z*�E]諽pb��UЩ�7B��T�
��St*n�MЩ�7B��T�
��St*n�M늽qW�*��^���z�\U늽qW�*��^���z�\Uޮ�qT�Q��S��*�W^��Z��늽qW�*��^���z�\U��σS��*��^���]w���uޮ���z��W]��]w���u-Wo����m���o\����-Wo�b�x6��m������σo��>�||�6��m������σo��>�||�6��m������σo��>�||�|�|�|�|�|�|�|�|�|�|�|�|�|�|�|�|��Z����Z����Z����Z����Z����Z����Z����Z��5�F���Q�#]Dk��u��5�F���Q�#]Dk��u��5�F���Q�#]Dk��u��5�F���Q�#]Dk��u���Q���Q���Q���Q���Q���Q���Q���Q���:2�v��]�-[��5�6J�N��W�h����59x�N^#S��Tp�*8hTQ��r��Q���[ b1�K$S�
=B�FJqJ�N)_)ǥ�LRE$ǰ$����JqIT�ϲC��P�)N�B��|vJR���W����~�^��߃¡�]-��bݬ6@q��n�?��G����3�E��n@~���M��O�Yt�՗O�Yt�՗O�Yt�՗O�1z������1 �?�l3��Ű�n-�+ql1[�}��_����~��+���.�$����S��Jw>N��)��hW>J?n�ܲC�b0���;J9҈�2#�IT���b��z�9���%�d�9C��(rx岾Q��Dh6$�Q��j1��&Z��J5Ij��Z����媟�j��Z����|�b�x1_>��������>��������>����-Ez�Q^��W��q���pk��?]���q���pk����q���pk��Ǯ[���p<o�[�����V��տ��o�-[��V��տ��o�-[��V��տ��o���������~}u?>���]OϮ���S����+�e�$F=�D�TN�w�NC��������m�x6��o�[�����e�2տ��o�-Kp�Է	-Kp�Է	-Kp��|'��	޷�w���|'z�	޷�w���|'����]�����~��}u߾���]w�N���]�Ӯ�t"�z_����N�S��Wbz؞�V3���Ec=u8�\V����Ei:ZN�V����Ei:ZN�V�����czu�ބV����T�{�;�NǽS����x5;NǃS����x5;NǃS���6�F�Z��KU	j�a-Tl%����Q���k�4���A���k�4���A���k�4���A���k�4���A���ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��$��d��l���]�O�I�v�?��'��$��d��l���]�O�I�v�?��'�P�;�;�ýC���oUu᷼5�N�>�Uӊ�7z��W]諽w���U���1W�*�T�
��St*n�MЩ�7B��T�
��St*n�MЩ�7�*��^���z�\U늽qW�*��^���z�\U늽qTJt�z���^���J4�e_\U늽qW�*��^���z�\U-To��n�js���ޖ�{�]w��uޮ�5�z���\�]pk�\����|娪Q�ݎTo������6��k��|�o��>�||�6��m������σo��>�||�6��m������σo��9j�9j���󖫩j�9j���󖫩j�9j���󖫩j�9j���󖫩j����j����j����j����j����j����j����j�����u��5�F���Q�#]Dk��u��5�F���Q�#]Dk��u��5�F*��Q�#]Db��u��5�F*��Q�#]Db��U(���Q���Q���Q���Q���Q���Q���Q��5�ʝj�vZ�ݔk�l�2M�7~)�#S�����5<6J��%F�F���A���P��(7��r��#��E"hQ��R�S�W�q�d��P��)^)�)�0e8����P��T(~��sՔ�z�/��O�I�m�u-�^�ߥ�w��f��v��g��h�[������g�N�}�����7O�$>��z*�B諉��$.����q!t_�B@W�E��$q(H
�P�X���e�VYH2�d1 Ű�o���J�h�3������^�@�`�	&�ip�'��I���|4(~��ߡC����$?v9 ׎C����(�"9�J1L	F)��Y�6�F�,���Q��9C��-���F�a���5�F�(�be��Q��j0R�O��Q��j0��O�S������|�b�x1_>��������>��������2�ẈS����2�W��]���n86�����׃]�����k�^v�o������~x2ߞ��Z�������F�	(�a%��j��Z�������j��Z�����b�����\V�S���z�~}qXO]O�J��E`c�8�NI)�,#��.�w�����]�-W`e��j��Z�������j��Z������nZ��%�nZ��%�n�o��[�;��N���o��[�;��N���o���~��}u߾���]w﮻��]�����a:u�N�W�B+���ީ�w�p]�B�ފ�w����g�����ⴜ��B+IЊ�t"���'B+IЊ�t"���'B+IЊ�t"��ꝏz�cީ���6����c����jv<���c����jv<���Q���6�F�Z��KU	j�a-Tl=u��A���k�4���A���k�4���A���k�4���A���k�4�j�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��r]�O�I�v�?��'��$��d��l���]�O�I�v�?��'��$��d��l���~�ýC��P�;�;�Uӊ�qWN*��]8��w��]M멽u7����ij���ij���޺��Sz�o]M멽u7����޺��Sz�o]M멽u7����ij���ij���ij���ij���ij���ij���ij���ij��@%���jZ<2�Q��+���T�e����\��Qpj.E���5�SKU4�KU4�KU4�KU4�KU4�KU4�KU4�J1TF�8�Fqʜ�4�J1T�J1T�]KUԵ]KUԵ]KUԵ]KUԣJ1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1TF���Q�#]Dk��u��5�F���Q�#]Dk��u��5�F���Q���
�|�A�߶K�1�6H��Y�"��Egd�����+;$VvJ��QY*k%Ed������TVJ��QY*k%Ed������TVJ��QJu5���TVJ��QY*(�M���9�*s��o��o�Tj�(7c�:1ʍ��X�F�F�V�A��Pp�(8b4q;%�����A��\P�}b4>�+d$F=	�}�G��QH�N)B�X�qJ�z�#��#�h�RE)�0e8~D�ȡC��;���sג~;%�)^�ߥ����=�_�~
�ip�^�@�x�x��X�}��?�[�a�܀�St�՗O�Yb̏��X��d��s��-�r�fK�QfK�QfK�]����+��\�Y�r�+���J@W)\d��ԥ��p�1!Ht����g�e�?���$?�[��Չ��Ŵ��[����q���+��M.$�v��ϒS��I0�)N�)��hP�YN�B�dP�H����Db�(���g�ȣ�9<r�'�hv�F�a��G(1��lr�(�c%Lr����*1��F
Q��J5)j��Z����a;��=�^ẈQ��j0���NC������|�b����V�����pb�x1XNW�+	�����a81_<�'+	���pb���'+	���pb���'+	�������1XNV����e���j��Z�����R�O����e���S�-E`����j+-T��QX)j��Z��KU?��V
Z�����R�V
Z��KQX)j+-E`�5߼��w����]������~�k�}qXO\V�]�����~��}u߾���]�'�o����x5��v2Z���QX�j+���*q�
�oB�Щ��*q�
�oB�Щ��*q�
�oB�Щ��*q�
�oB�Њ�t"���'B+IЊ�t"���'B+I����h5��_����h5��_��z�6�����a��z�6�����a����h5��_����h5��_����gz�,�Pe����C�z�ro]M-G���������r�z�Z�Y�Q�9j=g�Y�#�q���r=g�Y�#�q���r=gB�`Y q���Q�K84;ÃC����%d�Q�K%d�Z�����A���k�4�j�'��ryj�'��ryj�'��ryj�'��r~�ýC��P�;�;�Uӊ�qWN*��]8��w��]M멽u7����ij���ij���޺��Sz�o]M멽u7����޺��Sz�o]M멽u7����ij���ij���ij���ij���ij���ij���ij���ij����b�1	$��pj+$R��A�����nE���5���\��Qpj)F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b��Fq��4r��b�F*�b�F*���j����j����j����j��b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�b�F*��Q�#]Dk��u��5�F���Q�#]Dk��u��5�F��Egd��#]Y"��T�h4ezXf=����+;$VvH��Y�"��Egd��T
��PT*
�AP�*B��T
��PT*
�AP�*B���
I���
I��T
��PT*
9SG*h�Nq���%F���V�Q��݈�n�h7b4�J���/����Y(y��vJ�
��#C����P��(�6ϱg�%�&���⑲�R�S�W�qJ�MB�I��:;I����RMKVI�ג~;$���_㋿R�J�~N�/�K��v��_k�������Ϻ�������7O�Yz*�B�2?qYB,�yJ�9(�+1bVb<i��v�,J��X��ر+3�bVgbĬ�ŉY��2_Md��,�}7E��:)%i��J,��E��!o�P��ąV^��z-�;O�V$�� 6��gkm����.�$���J$�v�?�ϒI��I0�)N�B�vI0�YN�B�dP�H����P��6Kf��g�ȣ�9<r�'�P���F�a��G(1��lr�(�c"4؍69Q��Tc%��Q��j0R�F
Z����e���j��Z����媟�j��Z����e���j��Z����e���j������a81XNV����a81XNV����a81XNV����a81XNV�]�����a81XNVZ����e���j+-E`��������R�V
Z��KQX)j+-E`��������R�V
Z��KQX)j+-E`��������R�V
Z��KQX)j+-E`��������R�V
Z��KQX.O�������`�1X.V����`�v��]�'�]���c%��l��������'��Щ��*q�
�oB�Щ��*q�
�oz�Iި�w�4��'z�Iި�w�4��'z�cީ���v=ꝏz�cީ���v=ꝏ�_����h5��_����h5��_����h5��_����h5��_����h5��_����h5�z�,�Pe����C�z�ro]M��H�6������r�z�Z�Y�Q�9j=g-G����r=g�Y�#�q���r=g�Y�#�q���
�d�Y�#�iF�,������a-[+�d�Q�K%d�Q�K%��Z���4��Z����Z����Z����Z�����l���+�v��]���t⮜Uӊ�qWN*�E]��Sz�o]M멥��Z����Z��5���\��Qpj.E���5���\��Qpj.E����Q���Q���Q���Q���Q���Q���Q���Q�����W���ET(��A�z*�a��u7����޺��Sz�o]M멣�4r��T�ʚ9SG*h�M���Q���Q���Q���Q��5�j3�T�ʚQ���Q���Z����Z����Z����Z����Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q���Q������+;$VvH��Y�"��Egd�����+;$VvH��Y�"��Egd���SY*k%Md��U�t�{e�z����T�J��SY*k%Md���5
��PT*
�AP�*B��T
��PT*
�AP�*B��T�AI4
��PT*
�AP�3�Tg��������d�ղTj�j5l�x�풇F�A��Pe�T<4*�Ւ���C��P�"4>�[%�����C�B�BY#�VKdM
=)�#hQKNa$�$�LO$���{��s�J�MKVW�������>�Rݕ�8����W���;^����o!�!�����G�u:-�+z}q ſ�,��$->G�]+��2^J���V,J�G�#��6)��L�p��9R�r���@^�xT�6P��E�SY1Mg�#�>4��ŉY���Κ�|D-�r��G��q)B��B�?�/ESt�uo��S�-�:-�V!�����ez]��J�/�&��$Ըe?����r�n{��?vI�j�0�YN�)�4�P�"��Dc�6Ke���g�Ȣ6�dr�'�P��J|F�a��G(1��lr����h1�lr���G*1��F
Q��G(11dF�(�`�1_<����
=-T��U?��O�S�-T��U?��O�S�-T��U?��O�S�-T��U?��O�S�-T��U?��O�S�-T��U?��O�S����pb���'+	-T��U?��F
Q��J58�F+(�ce�l���b���V6Q���1X�F+(�ce�l���b���V6Q���58�F�(��e�L�S��jq2�N&Q���QX)j+-E`��������R�V
Z��pb�\�+���pb�\�+���pk���g�-Ece��$�S��jv<���Iި�w�4��'z�Iި�w�4��'z�Iި�w�4��'z�Iި�w�4��'z�cީ���v=ꝏz�cީ���v=ꝏ�_����h5��_����h5��,��e���A�ph2�Y���84d�C�KT94�C�KT94�C�KT94�C�KT97z�,�Pe����C�pm�.�E��H�6������r�z�Z�Y�Q�9j=g-G�����l�����z�Z�Y�Q�9j=g-G����F��Y�QI7=,��$��d��l���+娤�Z�Y�Q�>�E��H�t97��&����d��l�pm�.�E��H�6��"�ǥ��e��_�W���
��St*n�MЩ�7����޺��Sz�o]M-T��M-T��M���5���\��Qpj.E���5���\��Qpj.E(�R�E(�R�E(�R�E(�R�E(�R�E(�R�E(�R�E(�R�E)ð�c�{�WB��E^m܎�T�����޺��Sz�o]M멽u4r��T�ʚ9SG*h�M���4�J1T�J1T�J1T�J1TF�8�Fqʚ9SJ1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�J1T�Y"��Egd�����+;$VvH��Y�"��Egd�����+;$VvH��YЪ3�Tgd���5
�9N�|�C�+�(Ъ3�TgB�΅Q�
�:Ft*��T
��PT*
�AP�*B��T
��PT*
�AP�*B��T�AI4
��PT*
�AP�3�Tg����d�ݲPnШ2�*���/d��ШxhVʴ*�l�)��Э�(V�����l�d�@У�hV�J�S�}���T(�e
=)�#d�$���a��:Y+å���W��I79T��$Ե{����v��w�W(f�ߥ�C;]�����?$������u�-�+z}q �R>�qY��e��!ns����V,J�G�#��8�T.S \�@�WH㶝#��t�;i ^>�@�}��q��2�lj����@��B�9P�x�;-dv[ƕ��K�<i/������b��-�$(���z(b��C���H�:-�V!���-��a�]��J�~�'�~I�m��;��s����%x~��Ւaڲ�;>S�gРH��S�J�Q�%���l���%�d��C��P��:���#C����,�:K%��C���cb4��F29A��Pbc���2#C��j0^�������⑲�F
Q��J5)F�(�`���Q��j0R�O�S�-T��U?��O�S�-T��U?��O�S�-T��U?��O�S�-T��U?��$�S�-T��U?��F
Q��J5(�F29S��T�#�:H�N�9S��T�#�:H�N�9S��T�#�:H�N�9S��T�#�:H�N�9Q��Tc#���F29Q��Tc#���F2Q���58�F�(��e�L�S��jq2�N&Z���U8�j�-T�e��L�S���q2�N&Z���QX�j+(��%���S��Tl%����Iި�w�4��'z�Iި�w�4��'��c����6>����c����6>����a��z�6�����a��z�6����_����h5��_����h5�|�C�KT94�C�KT94�C�KT94�C�KT94�C�KT94�C�KT94�C�KT94�C�KT97��&����d��l�pm�)j=g-G�������b��SQ�`J1L	F)�(�0%����c�2�SQ�`J1L	F)�(�0%�F��Y�QI7=,��$������QI4���b��z�Z�Y�Q�>�E��H�6������r�z�Z�Y�Q�9j=g-G����=,�Ǥ������*n�MЩ�7B��T޺��Spj.E���5�QJ5�QJ5���\��Qpj.E���5���\��Qpj.E���5�QJ5�QJ5�QJ5�QJ5�QJ5�QJ5�QJ5�QJ5�A��)V#�ӷ�ԧ�$��t+�]M멽u7����޺��Sz�h�M���4r��T�ʚ9SG*h�M���4r��T�ʚ9SG*h�Fq��4r��b�F*�b�F*�b�F*�b�F*�b�F*�b�F*�T���9S�r�8�Nqʜ�9�*s�T���9S�r�8�Nqʜ�9�*s�T�ʚ9SG*h�M���4r��T�ʚ9SG*h�M���4r��Egd�����+;$VvH��Y�"��Egd�����+;$VvH��Y�"���7Ш*d���
���i&�:B��T
��PT*
�AP�)N���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN�|�A��A��A��A�d�ݡPe�T{%^�C�B�ڡP��v�R��ԧl�$ǱУ٨Q�Ҝ{���$Ǡd����S�}���RLR&I�D�1H�N)$�)$���������>M$���}����a��?"I���?�K������;��N�/~��żn���i��oE��b?k��Y�+}��ŜVB�YB,�yJ�9X�+14��x�;-qMMB�5����t�;i^>ǖ��>�5�"kzD,��Y���[ P�� P�� P��x�l㵵���^e�g�8�@\SYqML��oGi�.s�񳜔X��-�e�#�}q!HbA�ă��g�N�x�~������+Ըex?$�RےjW)_�I��Jw=yN�$õd�v�� Ҕ���(E�)*�G�(Q�$zMd�I�V�e
�'�P��:�%��C��P��:���#A����#���69A��h12�&Q���U.O���Q���m���Lr����(11�Lr����(12�F
Q��J5)F�(�`���Q��j0R�N&Q���58�F�(��e�L�S��jq2�V
Z��J58�F�(��c���F29Q��Tlc��F�9Q��Tlc��F�9Q��Tlc��F�9Q��Tlc��F�9Q��Pcc���69A��Pcc���69A��j1��F2Q��J5�F�(�c%�d�Q��j1��F2Q��J5�F�(�c%�$�S������N�Q��J5:H�F�9Q��Tl%|�Q���l=u]F��Q���l=u]FÃA���k�4���A���k�4���A���k�4���A���k�4��Z����Z����Z����Z����Q�H�d�Q�H�d�Q�H�d�Q�H�d�Z�ɥ��Z�ɥ��Z�ɥ��Z�ɥ���l�pm�.�E-G�������b��SQ�`J1L	F)�(�0%����b��SQ�`�1�F=�(ǰe����b��S9 ��b��RM��K81�d��KQI4� �G 2�SQ�`J1L	j=g-G�����"�b��SQ�`J1L	F)�(�0%�����$޸����z�n�Eި��z��T]ꋃQpj.E���5��j)F��j)F���3��3��3��3��3��3��3��3��3��3��3��3��3��3��3��3�Pg��9A�r�8�q���(3�Pg��9A�r�8�q���(3�I��(���ER�����t��gw�x5���\��Qpj.E(�Q��5�j3��g��#Q�F�8�Fqʚ9SG*h�M���4r��T���5�*h�M(�R�U(�R�U���4r��T�ʚ9SG*h�M��9S�r�8�Nqʜ�9�*s�T���9S�r�8�Nqʜ�9�*s�T����4r��T�ʚ9SG*h�M���4r��T�ʚ9SG*h�MB��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��I�NS��T���TT*
S��:�AP�*B��T
��PT*
S��:S��:S��:S��:S��:S��:S��:S��:S��:S��:S��)�o�Po�Po�P�ШthTyN���C�)�-Jt<r��l�$Ǳ�1�r�{D��$�.$��ē����x��&)$� ���L� �����R6I�RJ���^_߇����43s�J�<�������M�>W���?�K��܆`�p�׆-�v����B��t7��"����W����1g��l��ř/)E�Y%x�;MqLgd��H���@�}�x��5�e��j
�wj
�wzE@��K����*ˤT�H�.�P>R;�;�����;{ \��p;H�l���T,�P�MMB�55
Vi�.s�񳜔X��X��E\HZ�� ?Tض���:-�G�/�h���~�ߥ���~N�J�+�qJ�RO�d�ו���?^I�j�p��"I�dJqL%����Jq�4��P��z�OB�I�:��Od���(u�J|F�I��Dht�$r�(�be��r�d�RP��1�g��#C����"48ȍ2#C����"48ȍ29A��Pbc���&9A��Pbc���&9Q��Tc#���F29Q��Tc#���F2Q���58�F���G*1�lF����*61ʍ�r�c���*61ʍ�r�c���*61ʍ�r�c���*61ʍ�r�c���(1��lr����(1��lr����(1��lr����(1��lr����(1��lr����(1��lr�c���5:IF�I���*61|F�_���4���A���k�4���A���k�4�j�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryj�'��ryF�"�m�)F�"�m�)F�"�m�)F�"�m�)F�"�m�)F�"�m�)F�"�m�)F�"�m�)j=g-G�������b��S9 ��@0e����b��SQ�`J1L	F)�(�0%����c�2�{Q�`J1L	F)�(�0#�F)�-E$��RM-E$��RM(�$Q�u�r��`� 1����b��z�Z�Y�1L	F)�(�0%����b��SQ�`p`.E��H�0	z��T]ꋽQw�.�E���5�A��A��A��A�r�8�q���T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�T�(3�Pg��9A�r�8�q���(3�Pg��9A�r�8�q���0	x��&/B�Q�j(��4-�@�hw�hw�hw�hw�hw�hw�hw�hw�hw�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g���4�J1T�J1Tr��T�ʚ9SG*h�M���4F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�
�:Ft*��UЪ3�TgB�΅Q�
�:Ft*��UЪ3�TgB�΅Q��l��lP�*d��T
���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN���iN�|�A��A��A��A�d�ݡPe�:�
�jS���x�:i&ٚS�h��%8��&)q$�.$��į�+�?�0I&)$�"exd���`�L�I�RJ����:Y+å��|���E�<��U߹ʥ�)_�K��+Է{�}�f����$�~@o?"�4B@o(��{��qX�T�\V��s(E��P񳜔X���Gi�i������gΑ�ld����g P�[].��T�xڂ�
�����*������/P^&��MAx8���e�G���a�*˖���[��$
wzD,��.i \*�gʅ�e�.)��v�,J�D-�r�|���
�B��VY��Ű�n�[b��~-�E��xW~��ߥ���{��I�\����W�����;�=�^�+���v��ϔ���(t����G�(QI�=&�G��d��l�P����YB�K(V�=��_d���(u��F�I)�+��F�)�+��>���E,z�1�dr���G(q��dr���G(q��dr���G(q��dr���G(q��lr����(1��lr����(1��F2Q��J5�F����(1�$F�I��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a���*61ʍ�r�c���*61ʍ�r�c-P�e�l�C���q���Z���Tj�c-Ple���Q��h5��Q���(rx�O-P���O-P���O-P���O-P���O-P���O-P���O-P���O-P���O-P���M-P���M-P���M-P���M(�$R��E(�$R��E(�$R��E(�$R��E-G���������r�z�Z�Y�Q�9j=g��H�6��"��$\d��l�pm�.�E-[0%�f���c�2�{9�G"���RU�J��ITr)*�E%QȤ�9�G"���RU�J��ITr)*�E%QȤ�9�G 1����b��z�Z�Y�QI4� �G!�q~F*�åQ�r��`�1L	F)�(�0#��9 ��@0c��9 ��@0x0	"��$\��Qw�.�Eި��z���\�Z��Z��Z��Z��9A�r�8�q�������������������(3�Pg��9A�r�8�q���(3�Pg��9A�r�8�q��xv��Kjz�����VKe�j�������������������g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��9SG*iF*�b�F*�b��M���4r��T�ʚ9SG*h�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�:Ft*��UЪ3�TgB�΅Q�
�:Ft*��UЪ3�TgB�΅Q�
���Ӓm�N��PVJ��QP�)N���iN���iN���iN���iN��m�&ؒm�&ؒm�&ؒm�&ؒm�&ؒm�&ؒm�&ؒm�&ؒm��m��hwd���
�v�C�B�є�xe:ԧC�)���t<rM�D�l�)�4JqMLR�I�\J���S̯�+�?�1H)^+�#%xd� ��`�L�W�W�����:Y߇ɻ��43��nx0��D3s҆`���K��܆i|R����z-�l��~E�h���P4�t7��"����~��f���R>��J�J�9(�+14��x�;-qMMB�5���r�gP�}��B��-�}"�|�
l*
l �j4뗑�뗑�뗑����룦T/#i�GL�>^F�?F�.?'P^&�ƣ�xz��2�=�e�{d���.ix�B�5���ئwƑ�h�+1|�����諉O�Yd1 Ű�n@o)�n�?���.!��;���^�+��$���I�\��(g㋿s����L;VI�j�p)N�B�`У�(�
)"�G��H���l�P���N=&�[%�+d��l��(u�J}��_��C79��c���79B�vT/�d������6#l���#b6�؍�6#l���#b6���29C��P�#�8��29C��P�#�8��69A��Pcc���69A��Pcc��F�(�c%�dr����ht�$F�I��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a��Dh6�F�a(�)%e$�l��m����Q��J4;	F�a-Ple���A��h5��9C��(rx�O-P���O-P���O-P���O-P���O-P���O-P���O-P���O-P���O-P���M-P���M-P���M-P���M(�$R��E(�$R��E(�$R��E(�$R��E-G���������r�z�Z�Y�Q�9j=g��H�6��"��$\d��l�pm�.�E(ǰe����c�1Ȥ�9�G"���"9�G"���RU�J��ITr)*�E%QȤ�9�G"���RU�J��ITr)*�@0c�F)�(�0%��������iF"���"0��:U�J�0�Tr��`� 2�SQ�`G 1�r��`� 1�r��`�P�9jg-C��u�z��P]��Aw�.����4���\�AJ5�QJ5�Qph.���4���\�Az�)Fز@.�p��M�^���NZ���r��PQ�
9AG((���44F����#CDhh���44F����#CDhh������-��G���e8��z�%�vKd�4F���Q
#ADh(����r��TQʊ9QG*(�E���r��TQʊ9QG*(�E���r��TQʊ9QG*(�E���4r��T�ʚ9SG*h�M���4r��T�ʚ9SG*h�M��4F���Q
#ADh(���4F���Q
#ADh(���:S��:S��:S��:S��:S��:S��:S��:S��:S�%;bS�%;bS�%;bS�$��I�$��I�$��I�$��I�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$���&=VI�K�1�y^)�W�a��3w♥x��^=���ߊs��.!�Y^�W�u��exY^)� �$ÿ��ﲼ;� ��a���>�W�X����|����79d3�w��n�:���E�<g�"�ȋ~5bߍXf��  �R�� 6���_'~���t�t+O�Cb�t^@C����B�M���d�.,IyJ,IyJ�9_Gi�.)��.e^>ϤB�lt��2�=�����/PcQP|~N��:Νr�5A��ʇ��EC��"��l�Pr�H�~^�Pr�H�~^�Pr�H�~^�P\�2��<�q�7-�>[P6��d
�|�E@�rޗ{ P�[�|}�B�v���@\SSs��-�r��9�ř/%tX�����\[\H:}q ��:�Ca��6-�D!��*W���0~I&��$Զ��+�~�r��8����ݔ�R�J� Ȕ���?"I�J���I�J�8�� ���t(����Y#�k$zMd�I�6�dF='�Ǥ���#��c�x岾9��m�����Q�RDht�$F�I��Dht�$F�I��Y-�6Ke���cd�X�-�6Ke���cd�X�5�F����ht�Ke����`y&'���"4:H��#C����"4:H��#C��[+�9<r�'�P����9C��(rx�O�K"6�dF�,��%�d�#l�Dm�ȍ�Yd�K"1�<F='�Ǥ��e|r�_�W�4;岾9l��[+���岾9l��[+���F�a(��%��C��hv��Q���4�N�Q��Т�)&�+ò%8�F�"�j2�j�'��ryj�'��ryj�'��ryj�'��ryF�,�m��F�,�m��F�,�m��F�,�m���z�9��G���8�z�9��G���8�z�9��G���8�z�9��G���9F=�(ǰe����c�2�{Q�`�1�F=�(ǰe����c�2�{Q�`�1�F=�(ǰe����E%QȤ�9�D`Ȥ�9�G"���RU�J��ITr)*�E%R�S"Z�dKP	T� �KP	T� �KP	T� �KPj�-@0e�� ���2�Z�`�0�F�(ò%vD�Ȕa��;"Q�dKP	T� �KP	T� �KP	T� �KP	T� ����r�:�Z�Y�P�?]롽t7����޺Z���Z���Z���9AG((����Z���Z���Z���Z��u�CDb�С�e8}[$�r=9j��PQ�
9AG((����r����#CDhh���44F����#CDhh���44F����Kd�Q��Q��Q��Q����hh���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(�Fq��5�j3��g��#Q�F�8�Fq��5�j3��g��#Q�F�8���4F���Q
#ADh(���4F���Q
#ADh)N���iN���iN���iN���i&�9&�9&�9&�9&�9&�9&�9&ؔ�iNؔ�Nؔ�Nؔ�Nؒc�&<�c�&<�c�&<�c�&ؕ�ӕ�ӕ���������x��x��zr�z�^=9^=|����W�NW�_+ǯ�c�d��Y&=/+�0��L=���S7~)�W�h��9����Np��3 �+�:���2����߀��?��ﲼ;� ���0�>���w���}�~'�nr�f&�a�hf���!�~[s�C?oƬ[�Ի!����]������������� 7�?y��O�[b�q[��>�d�.,IyJ�9([��al��x�;-P��g-�v�"k`˥���(1��&����Atu�:��u%�Zu%�\�\��J�i�?�V���Zs��i�?�V���\�\۹b��iԖ���� ˣ�A�#t��PcQ�j��o-�}5����^e�g���B��M%f"�9X�%�>G��q!i�ă ?Tطy�w�طk@�v���/�W����~I&��Թ;�+����$��%x~���T(�|� Ҕ���;>I�J���S�`�p9NgB�H�QI
)"�G��H����Dm�ȌzO�I�1�<F='�Ǥ����r=c(�)%e$F�I��Dht�$F�I��Dht�%��cd�X�-�6Ke���cd�X�-�6Ke��Q��Pcc�؍������R�I�I�4:H��#C����"4:H��#C���l#�9<r�'�P����9C��(rx�O���6�dF�,��%�d�#l�Dm�ȍ�Y�K,�Ie�),�Ǥ���9l��[+���岾9l��[+���岾9l��[+���岾9l��[+���岾9l��[+�9<r�'��6����I0�	&*��1�9A�KT9<�C��T9<�C��T9<�C��T9<�C��6�d�l�J6�d�l�J6�d�l�J6�d�l�G#�q���r=g�Y�#�q���r=g�Y�b��F)��`Db��F)��`J1�F=�(ǰe����c�2�{Q�`�1�F=�(ǰe����c�2�{Q�`�1�F=�(ǰc�ITr)*�E%QDF��J��ITr)*�E%QȤ�9�G"���RU-E2%��D� �KP	T� �KP	T� �KP	T� ���2�Z�`�Pj�-@0e��Ȕa��;"Q�dJ0�F�(ò%vD� �KP	T� �KP	T� �KP	T� �KP	T� ����r�:�Z�Y��o]롽t7������-P��-P��-P��
9AG((�-P��-P��-P��-P��머4r=;$�v#�Q�%�#CDhh���44F����#CDhh���44F�����CY(k%d���5���P�J#AY(j�t+d�V�Э��P�
�CY(k%d���5���P�J#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
�CY(k%d���5���P�J�CY(k%d���5���P�JS��:S��:S��:S��:I�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�bI�$�c��ߊ]�Ǫ��{������z�~)w��ߊ]�Ǫ��{������z�~=VW�K��L2�S��ߊf��3J����>�S�~)�I�\J���S�~�� �߀��?���LW�}��=�tg~߇F����}�~'�����>M����?��C0���*�nr�sҋ~5dK^�vE�-ȶ����4��n���i��/�@q���{��|1X��wE#�g��ė��l�%%f#ƕ��Ge�.)��\Ӗ���2�����ڂ�
���0e��*��T<��i�snӟ�+�����n^+ d/S�2������rB�9!z����N�ȯI{-�s����T?��P�Z�Pr�H�>^F�&��H�	�(;�������/Ge�Ĭ���Y��9�W��rZ|���	e�k�������xgy��"��ߥ�J�~�^�Թ!��'�nW�ܥ8~�
�)�5�8�� Ҕ���;>� Ȓ`�&*��2�SS�`�qL{���G�,��5�=&�G��H����Y"�ȌzO�I���岾9l��[,l��%���l��[,l��%���l��[,l��%���l��[,l��%���l��Tlc����C��[$�zY)ǥ�LRMd���(u�J}��_d���(u�J}��_�K"6�dF�,��%�d�#l�Dm�ȍ�Yd�I���5�=&�G��H����Y#�k$zMd�K,�IdF='�Ǥ���9l��[+����zO�I�1�<F='�Ǥ���#��c�yj�_-[+�e|�l���ryj�'��ryj�'��k��#��C�T(t�� ��G��d�Q�H�d�Q�H�d�Q�H�d�Q�H�d�9��G���8�z�9��G���8�z�9��G���8�z�9��G���8�z�#���0"1L�S#���0"1L�SQ�`�1�F=�(ǰe����c�2�{Q�`�1�F=�(ǰe����c�2�{Q�J���Q�J��L��S"# ψ�3�0��># ψ�3�0��># ψ�3�0�F�(�3�|� ϔ`�>Q�dJ0�F�(ò%t�Q�J�t�Q�J�t�Q�J�vD�Ȕa��;"Q�dJ0�F�(ò%vD�Ȕa��;"Q�dJ0�F�(ò%�|�Z�ʥ�|�Z�ʽt7����޺�Cz�ij���ij���ij���h����r���ij���ij���ij���ij���\
Q�#���#ӎG�(����44F����#CDhh�d�N�l���;%�vKd���-��['B�N�l�
�:�t+d�V�Э��['��4���['B�N�CDh(�Ed���5���P�J�CY(k%��4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(���4F���Q
#ADh(�d���5���P�J�CY(k%d���5���P�J�CY(k%$�M�$�M�$�M�$�M�$�M�$�M�$�M�$�M�+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǯ�b���R^�K�1Ixf)/�%ᘤ�3��b���R^�K�1Ixf)/�%ᘤ�3���ex���~j�h�`;�N}��8fq�.%x^�:� �߀�aА�:�}�a�exw��>���ã!�}$3����!��|3s�C79d[s�E�93��nx2�"@|dH���� *Z�|v-�nH?3ې]�����q�"ݬ*-�´����G�/�:,���G�b�+!E�/)B��%�H�7�#����,�YP��-��pe=�l*������>^�P|�j��m?�+�wIA��2�I���3���;|�zv��������Cӷ·�o�{��8�I�q�;�Γ{�2B�>��[���-��J��ݧU�>��zeA��5A��82�r�����XYݨ^>���8�T,�Y�b�ر#�з9��X�KO���#�l1[�}�طy�w�طk@�v���/�W����{��K��rJ�;������L;�I�vI0�Y&�)ó�8v|� Ȓ`�&*�`�&*��2�SS�`У�(�
)"�E$T(����Y"��$RYd�K"1�<F='�Ǥ�J}��cd�X�-�6Ke���cd�X�-�4(��
=aB�XP��(��
=aB�XP���F�ad���(u�+d��l��q�d��Y(u�J}��_d���(u�J}��_d���#�k$zMd�I���5�=&�G��H����Y#�k$zMd�I���5�=&�G��H����Y"��$RYd�K"1�<F='�Ǥ��e|r�_d�K,�Ie�),�E%�H����Y"��$RY(Ǥ�zO(Ǥ�zO(�%���Y(�%���Y-P��Y�`Y 6H���`G#�q���r=g�Y�#�q���r=g�Y�#�q���r=g�Y�#�q���r=g�Y�#�q�F)��`Db��F)��`Db��F)��`Db��F)��`Db�Ȥ�9�G"���RU�J��ITr)*�E%QȤ�9�G"���RU�J��ITr)*�E%R�zU�dG"�ȦDF��g�`�|F��g�`�|F��g�`�|� ϔ`�>Q�g�0�F�(ò%vD�Ȕa��:U(åR�:U(åR�:U(åQ�~|r����!���~|r����!��;"Q�dJ0�F�(ò%vD�Ȕa��>U-C�R�>U-C�\c�lpm����86ģlJ6ģlJ6ģlJ6�F����#CJ6ģlJ6ģlJ6ģlJ6ģlph.-Pҍ�(���(�����44F����#CDhh�d�N�l���;%�vKd���-��['B�N�l�
�:�t+d�V�Э��['��4���['B�N�CDh(�Ed���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%$�M�$�M�$�M�$�M�+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧ+ǧߊ_ߊ_ߊ_ߊ_ߊ_ߊ_ߊ_ߊ]�`bإ��)j-�Z�b��إ��)j-�Z�b��إ��)j-�Z�b��إ��)j-�Z��3w♡��f�� �ù�0�fqàb�t~�� �á!�t$[��a�R�;�~߇Fw�ѐ�>���J���>���!���-�Ȣۜ���E�<��*�nr�?�WO�Ր-yR�����/sO�ܴ�]�@mw�.7�E��^�n�Ɔ��hoE����b��oE#�fG��ė��Ĭ��i����v⚙�6\���r�;{P��P^^��O,tu�:��j���U+c�%��u���K�]�2����Q�3�A�7�H�ä�a��0�~t0>� g�)�o�@�������"�u��c�!�Ǧ����~䊇��J���<�j*@�T.�� P�[ \vơq�/��B�S-ef#���V�#�z~+!H�6-�+l1X��������P%~4*�¡�_�~��p��6�{��I��Jp��N�$õd�v��Ք���;>S�g�0�&�$�2$�D� Ȓ`�SS�`�qL{S�YТ�*REB�H���5�=&�G����#��c�x�zO�I�1�<F='�Ǥ���#��c�x�zO�I�1�<F='�Ǥ���9l��Ǥ���#��c�x�zOd�K,�IdF='�Ǥ���#��c�x�zO�I�1�=
)"�E$T(����P��*REB�H�QI�=&�G��H����Y#�k$zMd�I���5
)"�E$VH����Y#�h��Y�K"6�e
)"�E$T(����P��*REB�H�QIr),�E%�Ȥ�9�G#�h�zM�I���4�l�G#�q�F)�d�`� 6HF)��`Db��F)��`Db��F)��`Db��F)��`Db��F)��`�c�1�F=��`�c�1�F=�d�J��IU�)*�E%VH����Y"��$RU�J���Z�J���Z�J���Z�J���Z�J���Z�J���Z�J���Z�J���9ȎE2#�L��># ψ�3��+$;J# ψ�3�0��># ψ�3�0��>Q�g�0�F�(�3�|� ϔa��;"Q�dJ0�F�(ò%t�Q�J�t�Q�J�����?>9ώC�����?>9ώC��vD�Ȕa��;"Q�dJ0�F�(ò%�|�Z�ʥ�|�Z�ʸ6����c�lpm�Fؔm�Fؔm�Fؔm����44F��m�Fؔm�Fؔm�Fؔm�Fؔm�Fؔm�Fؔm��zq���1K���-��['d�N�l���;%�vKd���-��['d�N�l���;%�vKd�V�Э��['B�N�l�
�:�t+d�4���['B�N�l�
�;%��V�Э��['B�N�l�
�:�t+d�5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d���5���P�J�CY(k%d��V�Э��['B�N�l�
�:�t+d�V�Э��['B�N�l�
�:�t(�I�$�bI�$�bI�$�bI�$�bW�NW�NW�NW�NW�NW�NW�NW�O����������������-�Q�a�b�u�F-�Q�a�b�u�V@@1�9 �  ���c�r�@@1�9 �  ���c�r��h�`!�����s�a�l;�[�àd?�3��aБl?�[����|~߇�C0��f��b۝�~a߇�E�h��M��R��-����T��ȐK_��k��~Ί���R�"�׋����[]�?k�w���E��1跑~�y�0Ŷ,���#�([%�qbK�^6s��vV�gj��k*q��/g�!f��g����C�8�X��=%+r�s+kZu%��\ҹb�������Qӷ·�h= o�����{�>��}��
��΅J@�B� s�RӷN��h=�� gr��P�N�v�v@�d���?��IjeAtu�[5����@�H,���Y��\v���5�bGi��s��YCO���>��t��A��t[V"�t^�C{�ȇy�v��f��Իa����ܯs�I7=�N�+��d�v��Ւaڲ�;>S�g����&�+ó�xv|�ϒ`LU$�%R�SS�`�p9Ng)�,�8�
)"�E$VH����Y"��$RYd�K,�Ie�),�E%�H����Dc�x�zO�I�1�<F='�Ǥ���#��"��$RYd�K,�IdF='�Ǥ���#��"��$RYd�K,�Ie�),�E%�H����P��*REB�H�QI
)"�E$T(����P��*REB�H�QI
)"�E$T(����P��*REB�H���5�=&�G��d�#l�P��*REB�H�QI
)"�E$T(����D`h�M�I�0	4F)"��$Q��#�Db��F)��`Db�H��B�J�1L�S#���0"1L�S#���0,�$� ��@0l�$� ��@0b1��{#��ǰb1��{#��ǰl�IU�)*�E%VH����Y"��$RU�J�0�F�(ò%vD�Ȕa��;"Q�dJ0�F�(ò%vD�Ȕa��;"Q�dG"�ȦDF��g�`�Hv���d�iY!�VHv���d�iY!�VHv���d�iG!�Q�v�r��iG!�Q�v�r����!���~|r����!��~Dr���G!���~|r����!���~|r����!���~|r����!���~|r����7<�F�(��%�G<�ǜ�pc�y(���(���(����"6�F؈���(���(���(���(���9J6ģlJ6�r<�@/�@/�G�H��Y#�$yd�,��<�E'B�N��
):Rt(��QIТ��ⓔⓔⓔⓔⓔⓔⓔ⓲[(�S�NS�NS�NS�N�Y-�yB�(Q�
<�G�(�P��%�d�,�Œز[Kb�lY-�%�d�,�Œز[Kb�lY-�%�d�,�Œز[Kb�lY-�%d���5���P�J�CY(k%d���5���P�J�CY(jyB�(Q�
<�G�(�P��yB�(Q�
<�G�(�P��^=9^(��^(��^(��^(��^(��^(��^(��^=8fv�Q�`a�fF�Q�`a����y���y���y���}>�O�s�����w=>�O�s�����w=>�O�s�����w=>�O�s�����w8f�-�s�a��w8��-�u�a�2����a�a�t$[����&@\�d�&���0��f��"۝�[s��nu��ξ@T�R��@\�d�@|dH��>���Գ��?f���{�/r,��P�k�x�1g���q�!o�!Q�[��şt~,����N��>��b���%�([��i����v@�L�p�[��D,���K��:��?/�g��nR@�-O�=s�3�o�?�+}G��:��:>�����j�P�s�P�s�Pܣ��nQ�T7(�*�w��;ʆ��|<|<���ā���@߆)�h=C�7�� g�+x^�����C�ܤq�9�2�����݃.�{�af��<��e�l��tY̥��yB@H�,[\H:}q[�a�Ā�#�o�/�!����aQn���;�~���ܯs�I0�)&�+��ex~�ՒaڲL?JS�g�p��N�߇�w��R�;>W�g����&�$�%RLU$�%RLU)�,�8�� ��E$T(����P�jMB�I�P	5
&�@$�(�� �Y"��$RYd�K,�Ie�),�E%�H����P�k$RYd�K,�Ie�),�Ǥ���#�РjMB�I�P	5
&�@$�(�� �Jp9N)�)�0e8�����2�SS�`У�(�
=�B�`P��(�
=�B�`P��*REB�H�QI�=&�G��d�#l�Jp9Ng)�,�8�� ���r��S�Y�`h�M�H�1IF)"��$Q��#�Y 1�F)��Y�b�H
�)ó�$� ��@0l�$� ��@0hP�U
*�C�T(t���P�Ҫ:UB�J��IU�)*�E%VH����Y"��$RUd�J��IU�)*�E%VH����Y"��$RU�J�0�F�(ò%vD�Ȕa��;"Q�dJ0�F�(ò%vD�Ȕa��;"Q�dG"�|F��g�!�VHv���B���!�VHv���d�iY!�VHv���d�iG!�R�;JQ�iJ0�)F�(ô�v��Ҕa��?>Q���0��F�(����D�sȎ\���=(��J9sҎ\���=(��J9sҔa��?>Q���0��F�(���~|�ϔny��"Q��J7<�j(���j(���j(����y�#��r<�G���9G#�$y�#��r<�G���9G#��y�"1I�b��G����"1I� С�l��<�G�H��Y#�$yd�(QIТ��E'B�N��
):Rt(��8��8��8��8��8��8��8��8��Q�
<�ⓒ`�0�8��P��yB�(Q�
<�G�(�P��yB�(Q�
<�G�(�P��yB�(Q�
<�G�(�P��yB�(Q�
<�G�(�P���t+d�V�Э��['B�N�l�
�:�t+d�V�У��t(�l�
<�G�(�I�(Q�lP��&ءG�M�B�$�b�I6�
<�m�&<��^(��^(��^(��^(��ӕ�^=9^=9^=9^=9^=9^=8fF�Q�`a�fF�Q�`a���Ԁ���y��7Es� .y��4��������d>㢇u�����@C�:(wY���d>㢇u�����@C�"��3��."�wX��-�@��f��BC0�H��-��H�L����|l3��a��>�-��ŷ;��c .u��ξ��$Ŝ����<?�U >24��~�R���Y�|�����T�ȳ�ⅻ]����<n?���q�:(b!Q�[��şt��G�o�d}6,g2�-�rQbVI^4���,�-P�O-�vU��A�K���PPcaP^'N�yNemj��w��t��{�2w(=&�Ǵ�Ѐr��A��v�Dw����(b@�� ~���?d���>@��G��H��/�Cqt��YGk�/�/�� o�sӷBN) gr�~�O����9�m�%�U��yl�H���/��*v@�f��q�(��jal��tR^J�YB@WE#�}q �_�v�V"�t^-�E���n���;�~�gㇿ�+��RL?�W�nJ���&�$õd�v��ϔ���;?��������)^�+ó�xv|� �I0	T� �I0	T����r��S�YТ�*REB�I�P	5
&�@$�(�� �P�jMd�K,�Ie�),�E%�H����Y"��$RYB�I�P	5
)"�E%�H��#��m�ȌzOB�H�P	5
)"�@$�(��� �P��*RE)�0e8�����2�SS�`�qLN)�B�`P��(�
=�B�`P��(�
=�)�,�QI
)"�E$VH����Y#�h��Y)�,�8�� ���r��S�Y�p9Ngd�Y� vH��gd�`� vH��d�`�b��r=g�`Y 4(D�ϲ@0l�$� ��@0l�$� ��C�T(t���P�Ҫ:UB�J�P�U
*�E%VH����Y"��$RUd�J��IU�)*�E%VH����Y"��$RUd�J��IU�)*��2%vD�Ȕa��;"Q�dJ0�F�(ò%vD�Ȕa��;"Q�dJ0�F��g�`�|F�d�iY!�T(~�
�d�iY!�VHv���d�iY!�VHv�r��iJ0�)F�(ô�v��Ҕa�R�;JQ���0��F�(���~|�ϔny��"9sҎ\���=(��J9sҎ\���=(��JQ���0��F�(���~|�ϔa��?>Q��J7<�F�(��%��������Q�%Q�%Q�"0F ��'�#��r<�m�Fؔm�j��G���9G#��y�#��r<�@(� P�
B�(P
 �@(� P�
B�(P
 �E'B�N��
):Rt(��P
 �@(� P�
B�(P
 �G�H��Y#�$yd�(Q�
<�[KbS��:S��:S��:�lY-�%�d�,�Œز[Kb�lY-�%�d�,�Œز[KbI�NI�NI�NI�NI�$�bI�$�bW�NW�NW�NW�%x��x�W�NW�$��I�;��w��&(�ǒLQ�'߇"����[ �~�`��'߀O�������]�`b�u�F-�U�a�b�uX�V-�U�a�b�uX�W��߇U�a���>^��ŷ<1l?[ǧ�h����r㞟��@|s�>���@C�d>O�y��>�@C�t�w�����d>O�y��>�@C�t�w���a�1l;�����a�a����-���a�d�&���78���I��"۝$������@\��ξ@\��߉<[�&�)����~,�۞��Ȑ}K?���E�?dY��tT��K����Z~׋������N�y��o;t��l��~i��EE��1m��;Ƒ�ر��=��Ŝ�P�vW��18�x��@�}�-�w������T?GYө-Zӟ�v@�L���/SӞ�F�����9}���<r��͒�?$����/ �+ &�dt��Rn�) ~�$�9�������������������r��H�x��ip��P���g�E9c�S�e�N|R,~�+r�#���/��^@��@�f����>[��.)���d~J,H�\-�,�c� şuo��[d/ 8�ދy������E���3�w������nW�ܥ�)&�$��;�=�^�+���x~�~�߇j���]�~�~�߇�w��]�~�� �I0	T� �I0	T� �I0	T� �I0�	N"���)N"���)N"���)N"���)N"���)N"���)N"���)N"���)Ng)�,�8�� ���2��S�`�p9N)�)�,�8�� ���2��S�`�qLN)�)�0e8�����2�SS�`�qLN)�)�0e8�����2�SS�`�qL$� ��@0l�$� ��@0l�$� ��@0l�$� ��@0l�$� ��@0l�$RUd�`�"��$RUB�dP�(E
�B�dP�(E
�B�dP�(E
�B�dP�(E
�)ó�8v|�ϔ���;>S�g�p��N�B�dP�(E
�B�dP�(E
�B�dP�(E
�B�dP�(E
��dD`DF��dD`DF��dD`DF��dD`DF����!���~|r����!���~|r���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F����!���~|r����!���~|r���DnzQ��F���DnzQ��F����!���~|r�(�'(��r�(�'(�'(�'(�'(��(��(��(���N#�r<�G���Q�%bQ�#��r<�G���9G#��y�(P
 �@(� P�
B�(P
 �@(� P�
B�(QIТ��E'B�N��
):B�(P
 �@(� P�
B�,��<�G�H��Y#�yB�(Q�
<�m�&ؒm�&ؒm�&ءG�(�P��yB�(Q�
<�G�(�P��yB�(Q�
<�m��m��m��m��m�&ؒm�&ؕ�ӕ�ӕ�^(��^(��^(�b�f(�b�f(�b�f(�b�f(�`� �`� �`� �`�>�R��R��R�fv�]�a�b�uX�V-�U�a�b�uX�V-�a�`b��������|�3��nxb۞��@\�H�r㜀���>���@\��78f������?�}���s������?�}���s� !�d?̀����2�@C���� !�d?�3���Ű��l?쀹���L3s��nq1mΒ-��E�;�a�XC?�_ .u�,��rh��M *R)�g >,�۞[s��}K?���tP}(�������� ){�~׋��\���&���距��@o?4�t+O�Cb��?U�G���+ ��/e�}�,�2�X�2���E��-xUB��}"�w`������>^�P�Z��?�T��+|0�N�@��n��@ܵ�9���9����@M+���Rޟ�A���3} O����d��A����T7���P�~V@K+�0�x���%q�h�1�iky~��Ix`sܶi�/]�/e�N��uC�4�2��u%�<���@Z�򀰳� P�[ \v�⚘����+%x�?%k�\X�H0���[�v����4_��E��47O�Cb�\B�»�/�g����w)^�r��8����~�߹�J��y^�߇j��ڽ�~�~�߇�w��]�~�~�$�%RLU$�%RLU$�%RLU$�%RLU)�,�8t�S�H�8t�S�H�8t�S�H�8t�S�H�8t�S�H�8t�S�H�8t�S�H�8�����2�SS�`�qLN)�)�0e8�� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	U
*�C�T(t���P�Ҫ:UB�J�P�U
*�C�T(t���P�Ҫ:UB�J�P�U
�B�dP�(E
�B�dP�(E
�B�dP�(E
�B�dP�(E
�B�dP�(E
�B�dP�(D�ϔ���;>S�g�p��N�)ó�8v|�ϔ���;>S�g�p��N�)ó�8v|�ϔ���;>S�g�p��N�)ó�8v}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv|r����!���~|r����!���~|F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��r����!���~|r����!���~|F���DnzQ��F���DnzQ��r����!���~|F �Ñ#D`��"0F ��# D`��N#�F ��# G"��Q�%�9G"��Q�#�Dr(�EȢ� P�
B�(P
 �@(� P�
B�(P
 �@(��
=}
=}
=}
):Rt(��QIР
B�(P
 �@(� Y#�$yd�,��<�G�(�P��yB�(Q�lI6ēlI6�
<�G�(�P��yB�(Q�
<�G�(�P��yB�(Q�lI6ēlI6ēlI6ēlI6įJ�D�J�D�J�D�J�D�J�D�J�D�J�D�J�D�J�D�J�D�J�D�J�D3 ��.�0���[�êŰ�/ !��/ !֤:Ԁ�Z��Rj@C�C0�xf/���۞��@\�E�=m�F����@��:�[��-���y�~<��?�|?���������|?���������|?���������|?������0�0�?�[���Ű��� .q2���"۝$[s��nv0�ń3�aԫ�ڕ~��'��rh��M�I�JE *R)�g�԰$Ī@|J���~�R���Qf�����:*^����]��q�Z~��o�[�س��衈�Y�P"��?U�[#�c�`.s!E��B��_s����b*�����q�)���2�=��j���<��9c��?�[�2����C���l�7���9-m`#�Cfe:�i_9����p�\�����|	�4��|��Ӻ@�l�������@�B�����Yj,��pşm?���-� %��g,�LV@咸���K�7z�TS��u=�]9�Hzu��*
V��%��#���/�P�_D�B�l�q���k<iY����1Y+��e[\H]1M��չ�����EƏ�\h��Ɔ��-��!�<*-�v�?=�����ܯ��+�qw�{����~��߹�C0�xf����~�3sՆnz���V������^�+ò%xvD�ȕ���;"W�dI0�	&�$ð$�v���a�L;I�`I0�	&�$ð$�v���a�L;I�`I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �I0	T� �P�Ҫ:UB�J�P�U
*�C�T(t���P�Ҫ:UB�J�P�U
*�C�T(t���P�(E
�B�dP�(E
�B�dJp��N�)ó�8v|�ϔ���;>S�g�!��Hv}��d�g�!��Hv}��d�gС�T(~�
�B��P��T(~�
�B��Y!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�!��Hv}��d�g�nzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DnzQ��F���DaȌ=�"0�F�Ñ# D`��"0F ����1I�!ӲC�d�N# D`��#�DF ��# D`��"0
 �@(� P�
B�(P
 �@(� P�
B�(QIУ�У�У�У�Т��E'B�N��
 �@(� P�
B�(P
):Rt(��QIТ��E')�')�'B�(Q�
<�G�M�$�M�$�(�P��yB�(Q�
<�G�(�P��yB�(Q�
<�G��zr�zr�zr�zr�zr�zr�zr�zr�Q+��Q+��Q+��Q+����	����'߀O� �~>�r�Q+��Q+��Q+��Q+���3 �èŰ�2/ !��/ !��}��sç�����z|?�ǧ�����ql?[s�����R�@\�H�r㞟���@��:�[��-���y�n�+�Es��p]����tW8.���\���>�O�����t��>�O�����b۟����-���8)s���"t���?�2-��H��a >,"ڕ|[R��jU��,��rm>�&�)��H��=�����X}K@|J���F�R���Qf��v��/v,�w4��Eƹt\k�Y�m�^���pşw�EB���Q�[��x�>�1Y�2B���#��%�/Gej��w*�q�.[6="�w`����?GY�>^FӪ���@�^��o��_R@�N,�ƀ��@M+�C2:Ԁ� ��\t��i� ]IܶKt�_�;��ӧ}A�4�?~��^�;���@�l����f�^����,�ʆ�,�+ %��Yb?����N��I�1�z�2{�%�T=sL�z�\�f@�����H�.�5��l�,��@\��I|���X���[\Yz(b������^�lY�[z-�_O�Cb�\B�¢ڗl[R�j\�����J�ߩ\���(g������"۟d[s�n}�mϲ-�׋~5�ߍx��_����������??����������?>I�`I0�	&�$ð$�v���a�L;I�`I0�	&�$ð$�v���a�L;I�J���I�J���I�J���I�J���W�dJ��^�+ò%xvD�ȕ���;"W�dJ��^�+ò%xvD�ȕ���;"W�dJ��^�+ò%xvD�ȕ���;"S��Jp��N�)��%8~D�Ȕ���?"S��Jp��N�)��%8~D�Ȕ���?"S�g�p��N�)ó�8v|�ϔ���;>I��I0�)&�$����~��Ғa�RL?J�ҡC��P�*?J�ҡC��P�*?J�ҡC��P�*?J�ҡC��P�*?J�ϲC����$;>�ϲC����$;>�ϲC����$;>�ϲC����$;>�ϲC����$;>�ϲC����$;>�ϲC����$;>�ϲC����$;>#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J#s҈���7=(��J��d�ղ|j�>5l��O�['ƭ��V#s҈���7=(��J�sY.k%�d���5��C�Hz���;$:vHt�����P��P��P����!ӈ�# D`��"0F ��# Y � � � � � � � � � � � � � � � �qK��R��)�.�qK��R� �S�_)�/���p�8�:r�:r�:r�:t(� P�
B�(P
 �@�Q)��Q)��Q)��Q+��Q)��Q)��Q)��Q)��Q)��Q)��Q)��Q)��Q)��Q)��Q)��Q)�LrLrLrLrLrLrLrLp��3 ��.�0���3 ��.�0��������������������������u^�:�3��a���:�[���Ű�ql?[���E���l?4[���E��r�@\�H�isͧ�s��9��:�ER��T��
��R� >!$�$������N����D��:�N����D��2� .pR� .pR� .pR� .pR� .pR���D����d����2��@|X��*�>�_�I�JY *R�R�H
��@T�Z|�O����,�����t�>�R����J,��z*^�EK݋;]ȳ����(��ۋ<nH[�ߋ0�Y�8z(b�C[������+�w�#�~4���)Y��)(@Y(@YY%@\S�x�WH��\�lzGK��/�P\~��%nSN��3N`�t�z�=���R>��,����uCrL��?�f�.;�h����<��
�Ӻ�:wT�N�:����.�Y;�d�H���P�N|='�׫N����P~.��D�5B��f�n>h� ��<�����I��fl��r�.@�z o��4Q�/d��Pm�N�rEAJ��x8��2�=�e��yo��X���J�4�q9�xج�$|�RESt�un,���V"����q��k@�iqf����!��$3R�j\�����J�ߩ\���(g㋿s����;�>��ϳ�s����;����y^�+��e�)_�JW�ҕ�4��)_�JW�����^�+��ex~�����2�?W�����^�+��ex~�����2�?S��Jp��N�)��%8~D�Ȕ���?"I���7<�&�$��䛞|�sϒny�M�>I���7<�&�$��䛞|�sϒny�M�>I���7<�&�$��䛞|�sϒny�M�>I���7<�&�$��䛞|�sϒny�M�>I���7<�&�$��䛞|�sϒny�M�>I��I0�)&�$����~��Ғa�RL?JW����=Y^�+��e{���sՕ�z���VS���w=YN�)��e;���sՔ�z���V�ҡC��P�*?J�ҡC��P�*?J�աC�hP�Z?V�աC�hP�Z?V�աC�hP�Z?V�աC�hP�Z?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V#Ո��b0�X�?V9ՎC�c��X�?V9ՎC�c��X�?V#s׈���7=x��^#s׈���7=x��^9ՎC�c��X�?V�sY.k%�d���5��C�Hz���;$:vHt�����;��N�v���������;$:vHt���!ӲC�d�N���;$:vH�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�R��)�.�qK��R��)�.�p�8��N|� �S�NS�NS�NS�NS�NS�NS�NS�NS�NS�NS�NS�NS�%8�S�%8�S�%8�W�%8�S�%8�S�%8�S�%8�S�%8�S�%8�S�%8�S�%8�S�%8�I�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�NI�_�.�0���3 ��(�0���3 �êŰ�1l:�[�êŰ�1l:�~V���0�xf/��Ű�r�@\�H�is� .y��D���=�@\�H��sѧ�h��4i�:*��ER��� t����jP�|O��i�/�}K�R��Ծ�U(Ί��T�:*�gER��Q�J3��Fi�:�N����D��:�N����D��:�N����D�U(ފ� >,t����R���V}J�����JY����|M����|�O����{>����A�b�.U�R�].U�A��(>|Y���ݮ�EK݋;]�[�ⅼn(��ۋ;͸[�ߋ��p��bT���E��~�ر\S�.+M񤽖�J�\�H�B�b�W�#���gzG���.�c�:]�H�ڃ�r�����KS9c�ӟ�~�ON�z>�>��j�,�Ɛ?)�x	����1g��,x�@^�@�W='T/�,@pf ��1�@�
��r�C8�x	��0t�d�1�h��3��A��P�N|='T��n���5�q��ρ4���9�Ҿs,G��K�9����l�?r��>)��qڃ��H2��|�j:D�t����>�@����j�+4���*s��YB�X���b��A���tY�+gym���?��Z[��E�XT[R�`��l~�rC0}��J�ԮQmJ��n�?����3��n�?��K��vJ�=Y^�+�iJ�R�Ɣ��+�iJ�]����s�w�r���U߹ʻ�9W~�*���]����s�w�r���U߹ʻ�9W~�*���RM�>I���7<�&�$��䛞|�sϒny�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R�Ɣ��+�iJ�R��VW����=Y^�+��e{���sՕ�z���VW����=Y^�+��e{���sՕ�z���VS���w=YN�)��e;���sՔ�z���VS���w=YN�)��e;���sՔ�z�(~�
�B��С��(~�
�B��С��(~�
�B��С��(~�
�B��С��~�F����a��~�F����a��~�F����a��~�F����a��K����d���.z�K����d���.z�~�F����a��~�F����a��~�F����a��~�F����a��~�F����a��~�F����a����F����nz���F����nz���F����nz���F����nz���F����nz�*��RP�/��B�P�j�B��B��B�]�C�С�hP�4(u:��v�s�d�ݲ\��a��a��!ӎC��N9�r8�:q�t���!ӎC�B�]�C�С�hP�(u�:�
v��B�]�C�С�hP�(u�:�
v��$�(�0	y&/$�%��� �$�(�0
2L�� �$î�0�L:��$î�0�Ht���!ӲC�)ç)ç)ç)çB�(P�JqD�JqD�JqD�P�
B�(P
 �@(� P�
B�(P
 �@(I�NI�NI�NI�NI�NI�NI�NI�NW�_+ï���exu�^vW�]���exu��:�~W� �߇U��0���{�=�uXfj���0�P�>^�Z�a���:�3�íC7<p��3s���E�=m�D��� >9��r��@\���Ys� .}d�=?㞟��@|s��W�ER��|�?�T�����tPx.���T�:*�gER��Q�J7��F�U(ފ��T�z*�oER��Q�J7��F�U(ފ��T�z*�oER���#4��Ί��T�dŎ�R���V}Jâ���(<�@T���,���m>&�x/O���T����A�z*\���ʺ(>|Y��E�^�Y�����^�k�v�����x�Qcyr���H[�����fᅰ�*,~�g�@���6,��𶸶řN���oƒ�X��PGd�,��@\S�xdx���u�e��`���T?�Ӯ^F�柧0m�����;��8||=Cr��͒�7�pş@��:N�[���Ӻ��zw��B�I��9e��$@K��ǀ�,@DA��RZp��x3PN��Y>�Yex�v�A��?�N�X�� ���@�B��x�cN?��7�Ju���>N��T=9��u۪
KV�˗��PcQ^����>[��*)����v�J�7���ė��̏��UąR-�S�o�a��E��[ȼ���$ց�aP�/���E�}������>�3ۆ`�qmKr-�nE�-ȶ��Է"ږ�[R܋j[���~�ƿ�_�������k��Z����3s҆nzP��J��C7=(f�������3s҆nzP��J��C7=(f��������sՕ�z���VW����=Y^�+��e{���sՕ�z���VW����=Y^�+��e{���sՕ�z���VW����=Y^�+��e{���sՕ�z���VW����=Y^�+��e{���sՔ�z���VS���w=YN�)��e;���sՔ�z���VS���w=YN�)��e;���sՔ�z���VS���w=YN�)��e;����$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ�sՔ�z���VS���w=YN�)��e;��
�B��С��(~�
�B��С��(~�
�B��С��(~�
�B��С��(~�F����a��~�F����a��~�F����a��~�F����a��~�F����nz���F����nz���r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�F����nz���F����nz��������d��|vY>;,��O��'�dF����nz����B�P�/��B��W5
�C�C�C�С�hP�4(u:�
F��V��F�s�d�ݲ\��a��a��a��!ӎC��N9�r8�:q�t��С�hP�(u�:�
v��B�]�C�С�hP�(u�:�
v��B�]�C��0	y&/$�%��� ��`�L�� �$�(�0
2L���$î�0�L:��d�N���;$:r�:r�:r�:r�:t(� JqD�JqD�JqD�P�
B�(P
 �@(� P�
B�(P
 �@(� I0	�0	�0	�0	�0	�0	�0	�0	����xu�:��+î��벼:� �߀a��0��{�=��~�� ���Ű�ql?[���Ű�ql?[����7<p��[s���E�=㜀�� >9��Ys� .}dϬ����>���O����9��+�?���y�^z/������A�(<ER��Q�J3��FtU(Ί��T�z*�oER��Q�J7��F�U(ފ��T�z*�oER��Q�J7��F�U(�?�3��F�U(ފ��Ԭ4����R����O�A���,���m>&�r.����R�:*^EK���1f�*�r���*�4�(�Kҋ4�X�K�趺�g��v�����7�(��B�w$-�rE�c���al1
�?��-�!����ş�~,���qX���oƒ�X��^4���,���q��w*��fΡ����v��� ���A��7,~㼱�����?�� o�s��Z��7�T7d���t^?,�c��;��n��ŧuC���ӟ^��&��0�7�@�n,i��?�t���PzqzN��;��"@�C�3�7P &�-80x�*��`%�r�=;��-t��^�;����w-�ܳE���[�T7$�x	b>�孬����@�TS�=�:���u\��ˣ�r�?�`ƣ����B��B�v��T,SSP�fv�8����P��"̏��UąR-�S��1X��ދy������E���3K��i�������_$3ۆ`�p�n-�\�ږ�[R܋j[�mKr-�nE�-ȶ�������k��5�����~�ƿ~��ߩj�7=(f�������3s҆nzP��J��C7=(f�������3s҆nzP��J��J�=Y^�+��e{���sՕ�z���VW����5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�?�OƼ��$�k�w=YN�)��e;���sՔ�z���VS���w=yN�)���;���sה�z��^S���w=yN�)���;���sה�z��^S���.z�K����d���.z�K����d���.z�K����d���.z�K����d���nz���F����nz���F����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����nz���F����nz���F����>;,��O��'�e�����d��|vDnz���F����0�����wЪW�nh�:q}�/�6K�%΍�V�s��C�Jw<r�����V�s�d�Ѳ\��a�b0��}��:��:��:��:��:��:��:��:��:�:�
F��B�Q�C�С�hP�4(uNVS�աC�С�l��H�$�vS�a����v9^�W��a��8vN�� ��C�С�hP�4(u:�
F��$�Q��we;��N�v����I��$��a��0��8t�8t��8�S�%8�� P�
)ç)ç)ç$��a��"��q�d�����+��ŰyyN9N9N9N9N9N9N9N|� �I�]�a�d�^VW�U���{��~�>�
=FW�Z�nz"۞�f�����E�=�?43���E�=m�D��� >9��r㜀�� >9��Ys� .}dϬ����^z/�������E������|�?��:�ER��|�5(H�R���_t��س��0xس��0zM>I���4�=&����z�[���z�[���z�[���z�[���z�[���z�[���z�[���z�[�����|�O�Xi�+>�a�Ԭ"ڕ|[R��)d��K4�=����{=>�����t�>EK�tT�WEK�tT�TY��E�^�-���ݮ�Y�vE�7d-�qB�7-�qE���,�6���n�7�/v�Y�8ao�,��g����6,���x�>�1Yƒ�_VJPGd�)%T)����w������ڇ�ڇ�6��9bV�4��ZӘ6�x^��٧n�>@��,�ƀ�S�$��d�?��,x2�
��>��u:K� w�i^D��P��i��5P�q$A�'N�p`"�K>���$�E��L�Y`"t�ӵC9�uPϖj��g�-�g4X�;�9$��~����Hs�uB��f����[�@M)��}��[];t>:M�:M��Ͼ�Pu�>��zgH�q=#���ޗ� \v�@��B�5����;M%f",�y+��rQfG��mqe��,W��V:/u�O�G� 8��f����!��~������>�3R�`�r�  �r�ԮQmKr-�nC?����[R܋j[�lv-��Ű}ض���b�>��_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�Ƽ�R��]��K�W�vJ�.�^��+Ի%z�d�R��]��K�W�vJ�.�^��+Ի%z�d�Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��㲅��B��|vP�;(_�/���e㲅��B��|vP�;(_�/���e㲅��B��|vP�;(_�/���e��d���.z�K����d���.z�K��F����a��~�F����a��~�F����a��~�F����a��~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~�r����!���~��sՖ�z���VZ���W=Yj�-\�e�����(�k�?�Ƽ��(�k�?�Ƽ��(�k�?�Ƽ����Ul�;�}�K�&�-�h�]hW9z�^�s��C�Jw<r���s�)��Юr�/��/��K�%ΌFv#��݈���a�b0��}،>�Fv#��ݔ��e8}YNVS�Ք��e8}YNVS�Ք��e8}Z:�
F��B�Q�@.�"�e8�&�W�����{�9^�I�ڔ��hP	z^��B�Q�C�С�hP�4(uNFS�ݔ�whP��P��P��8t�8t�}�L>�&|��� ��JqE
 �@(� Jp��p��0��}�L>�$Q!�u
G���;��bI��Ԫ�p��p��p��p��p��p��p��p�8�L:� �+ê��겼;~k��߇c�ñŷ=����ù��R�S7~��s�a���}�[s� .}d�9s� >9��Ys� .}dϬ����>���@\�Ś�$Y�BE��$Y�BE��$Y�}�5/�f������T��_��J,ԡ"�J���tPx([K����H[K������c�R�z*]�E���z�[���z�[���z�[���z�[���z�[���z�[���z�[���z�[�����|�O�Xi�+>�a�Ԭ"ڕ|[R��)f��i�{=>g���4�^���r���*�r���*�;\��K҅�]X[�Յ�]X���<n�[�ⅼn(���E���,�6���o��oŘc�,�0���Q[\P"�q��ŷƑ���%�c�`.s!xҲR��;%P�I*�H�B�2�#��T,����aP\~��%nS�?q�X��}%��M�4�й����e����d|����,���xܼ2�iݧ^���H�����M�*���R]'����1P��	�H��Ӻ���];�d�:Ӻ@֜I��HӇN,���qjH���:@ʆpf���Cl�'��ON���A�)[�4X� �E�CrL��3�9e�x���]&�à����/]�ݻ�r�Α���#����Y�.[ Y�ơg��#��Ge��s��2^J�\�E������j��+��-�S�/u�O�G� 8�طk
�i��/���Ű}�����ᚗ&�K���|��  �qmKr-�nE�-ȶ��Է"ږ�[݋`��lv-��Ű}ض�Ի!��d3R�j]��K��vC5.�f�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_�������k��5�����~�ƿ�_��+Ի%z�d�R��]��K�W�vJ�.�^��+Ի%z�d�R��]��K�W�vJ�.�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��B��|vP�;(_�/���e㲅��B��|vP�;(_�/���e㲅��B��|vP�;(_�/���e㲅��d���.z�K����d���.z�K����d���.z�K����d���.z�K����d���.z�K����d���.z�K�������nz���F����nz���F����nz���F����nz���F����nz���F����nz���F����nz���F����nz���F�(�k�?�Ƽ��(�k�?�Ƽ��(�k�?�Ƽ��(�k�?�Ƽ��(�k�?�Ƽ����!����B�f�T�Jp}*�k'�:K5
���R�B��B��B��B��B�f��0�hW9z�^�s��C��!�l���H}[$>��V��d�ղC��!�l���Hv$;����d�a�C��!�l��6Hv$;����d�a��%�0	x�^S�Z�a�%x~n��G~�W��a��8�N�S�a���e8vN�S�a���e8}X�>�Fv��B�]�@/�@/�@/��'$î�0�L:� �S�_)�/�E'B�N��F);$�$�$�:�
v���$�4Y�\P��e���$��� �0��}�L:��$î�0�L�� �+ê���2�;~k��߇c�a���w8��  �t�<$[R��`�QLt(�iN���߹�w��a�����-�@ſbڔ[��-���y�~<ſbߏ1oǘ��ΟR��Ծ��/�}K�R���D��:}K�Y�BE��$Y�}��x.��A��6,��am.���z(=E���������Pz��K�Ś\�,���f�'�4�<Y����.Oirx�K�Ś\�,���f�'�4�<Y����.Oir~�_�A��(<�����O  �yR�H
��O����{9���x|��ʺ*\���ʢ��",�r"��",�r!n�V�uz-��Y�vB�7-�qt[�.�y�w�qgy�}ܐ���a��p�P�*,��g�@���6��[\[an+[�^��I{,X�d/VJPGd�)%H)��X���pJ��w��z4�e����̭�i�n�/e�@��N�8|��]K�YG�-�j��f�.:@�����*�N����ykN�;w�"�7P�����U�O����8�w�5 u w���C=8���8�I�8���8CU��rϧ@�MC
���N���i�;�M"܁@@�-�;��#@��I�"�:�q�p��t�̎�3)⼲�P�x�t�rz�������R�H�|�PcQ�:_mB���8��^eqMg�#�з9�E�/�褼��b��-�$([\Yb��A衊lY�+�ۧ�"���iqgk
�v��f���x{����/�Kߋi|�m/�-��C0}�f�����}��r��C4�(f������^�3K܆i{��/r�݆~7a���g�v�݆~7a���g�v�݆~7a���g�v�݆~7a���g�vI��~;$���'�I��~;$���'�W�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvS�n�u-�N��)Էe:��Rݔ�[��Kv���B��|vP�;(_�/���e㲅sܡ\�(W=��r�sܡ\�(W=��r�ݲC�l���$?v�ݲC�l���$?v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�vQ���7=�F�(��e��sݔn{���vQ���7=�F�(��e��sݔn{���vQ���7=�F�(��ex?�&��W���w�d��Ƅ�ôw���MJS��I0{�K��R�B�s��\�:�:K4�R�$�f��0�w<t+��
j�s��C�P�r�(}��^��B��С��P�T(}�>�
j��B�ڡC�P���P�VHv$;����d�a�C�P���P�rL;D��+��w�z;�=�?4��$ñ�p�2�;��)ð�p�2�;��)ð�a�b0��(u�$�$�$��Rq��x}^FI�]�a�e8��N|� �� �� �� �� ���B�]���e8}�Rp��[K�B�]�G�(u�NF� �W�ѕ�wex}^FW�ѕ��exuY^���߇c�ñ����w8f��s�a�a�����/���W�\I0}�X���3s��np0��-���y�~<�
��R� *_�K����/���@T��
��R��A�(<E���]J3��FtU(Ί�`�P�����.&,��b�.&��!m.�,ml"���,���f�'�4�<Y����.Yir�[��Bݬ��e��k,��Yd-��!n�Yv��[��Bݬ��e��k,��Yd-��!n�Yv�ȳK�Ś\�,��f�,��r�>�,���m>&�x/O��t[\��*�r���ȋ;\���ȋ;\�[�υ�l���׋mx���<n�[�ⅼn.�y�}�(��ۅ��H[�䅾�H[�텿�س��E��B�ر#��bG�"ď�E�/M�^�d��,g2��*��IR�ed�Hq��.cP��P��N�EC�u�:�ծ��d83�"�g�P��й��ip�!�3=�Vޟ�r�af��+zO�(^Ɯ� �iڅ�-ӃoN�"4",��$�Ĩe>�]8Y9gӁ��T5���*Ӂ�pi��q����@D����i�ӍP�C9R]'�D�E��N<X�g4X���,�P�@ܣ�}A�:O�Z@�-�f��i&V@KB��v����)pg�E9c�S�86�R��\}3�x5���y�����\�cP��W�#�1bVgb̗�tR^J�\�Y���[\Yb��A衊lY�+�ۧ�"�~�/�hnց�aQn��a��3��v�2k� 6��k���"�_$3ۆi|P�/���C4�(f������^�3K܆i{��/r-�nE�-ȶ��Է"ږ�[R܋j[�mKr�݆~7a���g�v�݆~7a���g�vI��~;$���'�I��~;$���'�W�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��Kw�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��rS�n�u-�N��)Էe:��Rݔ�[��Kv���B��|vP�;(_�/���e㲅sܡ\�(W=��r�sܡ\�(W=��r�sܡ\�(W=��r�sܡ\�(W=��r#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�v#s݈��b7=؍�vQ���7=�F�(��e��sݔn{���vQ���7=�F�(��e��sݔn{���vQ���7=�F�(��hP��O���J'�Ƥ��Ԓ�c =ђ�
W��J{_���
��I���R�%8=�
��S�s���%:�:K5�E
���s�d��d��|c�\�Y>1�.y���<�K�iN�S���y�;�iN�S���y�;�k$:Ւj��B��C��w<ҝ�4��I�h�����;����s����%x~i&�S�Z���8�NjS�a���e8vN����Q�è�a�l��H�$�vS�Ք��exuY&FI�Q�`e8��N)v� �d�]�C�С�hP�2�>���)��� d������d�]�C��p��(u��ί~�W��������~�>_��߇��ñ�0�p�;�3�úŰ�l;�[���{��f����àb۟���o)!�����-���n��$�����}K쀥����  �R  �R  �Z}.7O������>����t�\n���0xرK����[K����H[K��[����[[��Bݬ��dзk&��Y4-�ɺ-����ɡn�Mv�h[��Bݬ��dзk&��Y4-�ɡn�Mv�h[��Bݬ��dзk&��Y4-�ɢ�E8�(�ƑE�4�,�l����,�l���Ϣ���[\��*�r��Kҋ4�([�Յ�]X[�υ�l���׋mx��ׅ���[�݅���[��˔Y�mŝ��-�rB�w$-�rE�c~,W�g��?��-�(bG��lV?$}c��i�bK�|l�A�̅�J�\��*��IP�@\S;�xUAq�=:��:�~X��:��nX�i����J���$�� #�o %�H�	���7E����I�"Ӿ��PzM���,["�Hӏ�t0:pt�c�ā�Y������yR�r��',�p�dӍ�$��8Y9gӀ哖}8�P֜,�qj�cL�8d���6�H3r"XfD�����,z��T�w� ��\t��R:���Z�:M����4�Q�x6[�)-O�.�H�.>F�.�@�EB�6p8��,�qMdX��س%�+��2^J�2?$|�k�,Y�H:|1X��n���������Cd 8�	ƈE�nط���b�7n�������k� 6��k���"�_$[K�i|P�/���C4�(f������^�3Kܐ~)�~)�~)�~)�~7a���g�v�݆~7a���g�v�ݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݕ�[��KvW�n��-�^��+Էez��Rݒ`��LrI��I0}�&�$��$�>�ܒ`��LrI��I0}�&�$��$�>�ܒjW)&�r�jW)&�r�jW)&�r�jW)&�r�jW)&�r�jW)&�r�jW)&�r�jW)&�r��8�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S��\�(W=��r�sܡ\�(W=��r�sܲ|nY>7,��O��'���r��d�ܲ|nY>7,��O��'���r��d�܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��ܔn{���vQ���7=�F�(��e��sݔn{���vQ���7=ر#�!mq*�?���,�`�M.2�X�R>�������R�
I�BJ{_�-�Z׭��q)��$�=ē��`��K��R�)Թо4P�4P�4P�4P�4P�4P�4P�4P�4I?$��OƉ'�D��I��$�h�~4Y!֬��T(~:?�s�$�h��\�z�9&�W�����!�����^���W��a��v9&�I�c�a��}�&jI�ڒa��W9z�^��d�աC�С�hP�4(u&�/)����겼:�� �$�(�0
2�R�v��B�Q�C��p���>���$���8}YNVS�Ք��d�����)���p���|�~�W��������~�>_��߇c�a��w8��-�u�a�d?̀����2��~���0�0�?ΟR��o)9mq'�n�۟��	 >!4���>��O�}��_t�\N�����q:}.'O������>����t�\n�K���q�}.7O������>I���!m.����E���X��ō���ư���7�,q��c�&�iX�H��E8�(�ƑE�4�,q�Qc�"�iX�H��E8�(�ƑE�4�,q�Qc�"�iX�H��E8�(�ƑE�4���Y���?yg�o,�o�!o�:-�Y�J���",�r!n�V�uan�V�ub��J,o4��_��vB�wdX�7bǻr,{�"���7�(��ۅ��H[�䅾�H�oŘc�,~����B��$|7��c�K�|lV�d�o��d9�b�s!xҳdvJ�b�T�18�t�eP~>�N���<F��9=:��m9�m�s��J����ӷ��,G����M���K�uB��T��,x`"���"��[Pϖj��:�1�8�w�OP�N=C\��I�c�<�`'�k�z��r�Pԁ����j��������Y��r� k�NY*��N',�wT1�;��N?,�"]>D���]9��T�������B���q
K�C-~�M��t���/�N�6�2�����]#��t����^>¡gڅ�l�8��\SY%fZ�:h�%�fK�P��"ď��mqe�?���S��b��{��~�? 8��Ɔ������H���~H��[���ߚ~׷O�p��n�ߐ]��ߐ]��kr�v�(�kr�v�(�kr�v�(�k��x��]�O�ܴ�]�O�ܴ�]�O�ܴ�]�O�ܢږ�[R܋j[�mKr-�nE�-ȶ��Է%z��Rݕ�[��KvW�n��-�^��+Է{�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����;�}��s�����$�>�ܒ`��LrI��I0}�&�$��$�>�ܒ`��LrI��I0}�&�$��$���I�\����I�\����I�\����I�\����I�\����I�\����I�\����I�\����I�\����I�\����I�\����I�\�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S���8�?�)O�S���8���O��'���r��d�ܲ|nY>7,��O��'���r��d�ܲ|nY>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7%��sݔn{���vQ���7=�F�(��e��sݔn{���vZ�Fw��([#���q�+�e���%J�������%tl���h\hK&��Gkօ��$����2�̓R��jP2MJS��)�u��:�e?����YO㬧��S��)�u�~4I?$��OƉ'�D��I��$�h�C�Y!֨P�r��4��W�s���;�{�N�S�\I7;�_㬯��I��Jp�r�?�
���B��C�С��P�t(}�>ԧs�)��С��P�T(}�$;��)ð�0�RL>ԯ�+ð���2L^I�K�0	z^� ��@%�8vN�S�a�a���}�^玅 ��@%�}���i^�I�ڕ�0�7<0��3s����7<p��3���E�����-�@��� !К|?���������C0�Hf	 .pQckc PĲ@\��
@\����?�'O���Q����t[X΋k�mc:-�gE��趴�֓���t[ZN��c�R�z*]�EK��v=.�,mlb�����Xx�k�_w�x���]�,q��c�&�iX�H����,�l����,�l�m埍���~6����Y���?yg�o,�m埍���~6����Y���?yg�o,�/���"ǻ,{�"��,o0b��",o2"��",�r"��"��n�V,q����^,�5���K��j��wd-�vE�cv,C�cݹ�CQg�r�>�-�rB�w$-�rE�c~,{�b�1��W[\P"ď��ج^,b��K�`,���Y/[���d���^4���lRJ���V�gj��e�G��>;��Ö<GIq��X��N��ҺK�o�(^�TSN޸?,�t�L��? 3��c����z=;��c��zpd�:q$��`�P�,��	���E�jx����j�����OPʡ����OP˖z��r�Pԁ�Y��j�����j@��Y 'ӋP�L	���:ӻNt�T7t�����K�b��]'T._N�@M��г��K_���md�C�K�AӯM������z�q�ΑP122��oj�����,b��Gjans��2_d��qYB,H�
,H�
,��������E��^�n�����Ⱦ����O�P$! 7��y��q�:.7�E�������O�p������Ż[�[��E�[�[��E�[�[��E�[�[��E�[�[��E�[�[��E�[�[��E�[�[��w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�J��)^��+���z_�K��|R�/�W��J��)^��+���z_�K��|R�/�W��J�}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r�nW���p{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���P�\T*�
��B�qP�\T*�
��B�qY>7,��O��'���r��d�ܲ|nY>7,��O��'���r��d�ܲ|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎|nJ7=�F�(��e��sݔn{���vQ���7=�F�(��e���Jq؞}�~��%�t�V�+�����?����Wž�g���D��h)N�	)�Щ~ez\$�K�����?�^�S�y�j^e8<�R�)��d���N$Լ�px&��I�@�?$��OƉ'�D��I��$�h�\�,���j;D��$��;�(f������L?����W��+�u��:�7;�N΅�B��C�С��P�t(~:?
�I��$�h��y�;�j?
�I�c�a��v9&�S�Z���x�S��B�a�@%�P	z^S�a���8v&�I�c�~9Т�l��y^�-�\w�z%x~n��D��+�����Ҽ?4��+��J��r�?�~׿��a�a��f	��Ű��l?�Y�����ފ�߹���!;�?�fI=����Ai��mJ'O���xΊ�  �֓���t[ZN�k�mi:-�'E��趴�֓���tT���c�R�z*]�EK��v0��_x��7���.�O7�z���x��X�I��M8�(�ƑE���Y��ŝ��Y�����?yg�o,�m埍���~6����Y���?yg�o,�m埍���~6����Y�_vX�`E�vX�`E��X�`ō�DX�dE��DY��B�6|-�gŎ6�X�kŝ�Y�k���_ݫ}ݑb݋��X�7|hc�Ɔ8�Ϻ�}�([�䅾�H[����X�pŘc�Ʈ(bG�bď��ج_ƒ���� ,���Y/[��2X�e#�^6)%@\�+P��5B�2ܷ��T,�T?��Ӟ?�g�%nS���wI{-�s����ӷ��,G�,�%���o�@A�I�u�0�?CN��'N<��t��t����j&,��$�5�',���Ӏ�@֜,��� '�kN5C\�T2�@�C.Y9d�L��5 j}8���ƀ�N$����5:M"@���Y&�It��?gI��Ӈ���C<,�����Z�$�R��C����Ǌ�PU�*���>��g-�9��x��j�����,b��Gjans��2_d��qYC��qqbG�P����P�7O�V�/u���[t��_O�E��t7O�Ct��O�P$! 7��gy
�ߝ��~i�^�?�ç�d�~-��E�[�[��E�[�[��E�[�[��E�[���m�6܀�m�6܀�m�6܀�m�6�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�~�߃�w����>�K��|R�/�W��J��)^��+���z_�K��|R�/�W��J��)^��+���z_�ە��r�nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܧ�Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{���Jp{�
��B�qP�\T*�
��B�qP�\T*���r��d�ܲ|nY>7,��O��'���r��d�ܲ|nY>7,��K�s�r9��܎|nG>7#��ύ����s�r9��܎|nG>7#��ύ����s�r9��܎\����˟s�r9s�|nG.|Qύ��ϊ9���G>7#�>(���s�r9�-|nK_������܎|nJ7=�F�(��x7=��s�sܔa���?s�s����87=��s-���$9Jԏ�Xx����q
�g�+8����EƯ�4�H�d-�Xi����2W�D�5�����e8<L��F�>��O����K���p���K��jP�(?�&�	)��a�_YK��iw�=ē��jP2��Z��R�)Լ�?䟏�MK̓R����������ߩ@��P2��Y_㬯��I��I7;�N�S�����89N�S�����89&�q$��$��ēs��nwM��I��I7;�&�q$��$��ħ�+���p�rL;E
���B��C�С��P�(~:;E
���)���p�r�?��s��nwL?���$���0���?̯�+������?����^�s�߹�����?P��3�ԢdJ6�Fŷ:Hf� >,d.�,��������
]�E����_ )v=������zN�kI�R�z-�$Y��E���Y��B�5|Y��B�5|-�W��5|X�I���O7�x���Ŏ4�,�$�6�E}�/y"�Ŝ�`E�vX�`E�vX�`E�vX�`E�vX�`E�vX�`ō�X�`ō�X�`ō�X�`ō���x��W��x��W��x��W��x��W��E�bU!�TX�%Qb�E�bU=��cݟ=��cݟ=��cݟ7�Qcy�7�Qcy��o;<m�g���񷝐�y�w�����x�Qcyr�˔-�rB�w$-�oŏwX�pŘc�Ʈ(���E��>1X��%�KӢ�s[����s�ƕ����(�b*q��.;P�L�y\�����G��3�LӴ/n�7���^�UC���w(0�a�=py���r�+4[�r�<2+t�f��%Ӑ;�7B��P�-Ӊ {����E�?>�X�q�T1���=C�	<��1�~Y�$�O k�z��@O>�h	�Ӎ=CR�H�5�%C\�H���$�	j�ӏ�t0j�U$w�O�.I�܀� R��Y�`&�s��<V@ܣƀ����o:@���P�N���n���>��dq�5AA�ύ�wj���\���9^4�����Md�",�y*Ⲅ-������Qg��)M���E��t_�t��#����Ⱦ�����ȼ��Cd 7�?y@���	ƈH���~E�nط���a��3�߆v����~���;]�gk��w�_3K�i|P�/���C4�(f������_3K�i|P�/���C4�(f������_3K�i|P�/���C4�(f������_3K�i|P�/���C4�(f�����x>ܯە��r�nW����}�^�+���x>ܯە��r�nW����}�^�+�����N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����%x>ܯە��r�nW����}�^�+���^ܓKےi{rM/nI���4��&��$���^ܓKےi{rM/nI���4��&��$���_*�ʅ�r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�U.*K��R�T��U.*K���r�|\��>(���Q��z��?rS���t���ϊQ��z��������$�xhP~H����Rێ\���>(���#�r��\�~���k�_R���sۖ�8���ܵ��-\�寎)j�-|qKW=�k�Z���_R��nZ��|nK_�>�Kܖ�w.�9s���,�>)j�����{r�K~Z�o��/��s�����w=�]�o+�VP�e{>�(U�q1����3\rT
�>n@�]-?�,�jV=���Y�H���諉f����b�W��P�"h_=�������u(�N)��e:_����A��px����J����/�����^e?����O�����S����d���O���������~�ߩ@��e����Y&�q$��%89N�S�����89N�S�����Y&�I���a�d�Y&�I���a�d�Y&�I���a�e8uħ��@9Р�89N�S�����89N�S�����8uħ����L?���$�����2�?̧����>S��I7?�M���+�AI7?�M��s�+�AJ�R��~�ߩD��);����6W����)!��������Y<����
]|����
]|����
]|����
]EK��v=.�,�l"���,�l!o���o���o�,o$�cy'��?��x��d-�Y���-�Y���X�`E�v�`���X�`E�vX�`E�vX�`E�vX�`E�vX�`ō�X�`ō�X�`ō�X�`ō���x��W��x��W��x��W��x��TX�%Qb�E�bU!�TX�%Qb�E�v|X�g��Ɨ�ix�Ɨ�ix��_ݫ�{�|ov��n�_v��n�_v�X�nE�v�X�\�����{��ov�-�rB�w$X�pŏw�v���o�\P!mq@�>$|6,b��K�b�s[��n�2�d/VJPGd�.)��Yƚ@��B�s�c��xгc�<��IlN���GIzk\����?�;�o}F@�� o�R�7(�%�b��8�,�g��= \I���;N|5$� "�7�@H嚡��"���N,�Y 'Ӌ j~Y�'��x	�g�j~Y��5�=CU�g��N7,��2���~Y9d哖J�R��H��P�,�9gӉ������M Pf$E�'��N���� R��Y�`&�s�	d�/ nQ�iۃR�3��?���P�N��rAIj-��#����x�����.i�g�Ge�ns���_d��qYB�|\Y�d.�G�z)M���E��t_�t��#����Ⱦ�����ȼ��Cd 8��?y@���	ƈH4B@o?"�7l[��xݰ�׆���;]�gk��wᝮ�3�߆v��n���nQn���nQn���nQn���nP�/���C4�(f������_3K�i|P�/���C4�(f������_3K�i|P�/���C4�(f������_3K�i|R�nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��}�_'~��ߥ�w�|��_'~��ߥ�w�|��_'~��ߥ�w�|��_'~��ߥ�w�|��_'~��ߥ�w�|��_'~��ߥ�w�|��nW����}�^�+���x>ܯە��rM/nI���4��&��$���^ܓKےi{rM/nI���4��&��$���^ܓKےi{t/����B��P�.T/����B��P�.T/����B��P�.T/����B��P�.T*�
��B�qP�\T*�
��B��P�.R�?r�Rۈ�\�0�j�d�o�*[�}��R۔a���;v#�r�\��qM~�{VZ�n�`��;vZ�n�.|Q�����B��P�����nZ���W=�j�-\�嫞ܵsۖ�{r��nZ���W=�j�-\�嫞ܵsۖ�8��������v���/rZ�ܢ5.+%ϊ�v�;^j�йܼ1M�{r9�T�}w=����z��޹�J�Ku%k���#'PrW�zw>ȏs��y"Ďۋ��E�Ȇx�p��OB��J�h->���2>M�CqoMߥ�䚕���_$Ԭ,�*K$&#�����i~h[^��4$�K���p��.���A�(U(+'��J
�R��~ ���)^�	�BC5/��K���$Լ�5/2MĶ�)�@�4+�Zϭ
�օs�B���\�Ю}hW>�+�Z>���C�hP�>���C�hP�N��S���C�hP�$;�����d��Jp�r�?���)���p�r�?�������:�S�\I0�&+�����2�?̯�)��%8|$�s�$���7?�����+�AI7?�����+�Aw�Q=��O~�ߩD��);����6W����8���$[����?k'���}?k'���}?k'���}?k'���~��cv�gkav���_x��_x��_x��cy'��?��x��g��x��d-�Y���X�`E�vX�`x���`����`����`����`����`�����x���ݟ�{��ov������7�?��g����ݟ�{��ov������7�>,C��J��1*�Ī,{��ǻ>,{��ǻ?Ɔ4�hcK��j���_ݫ�{�|ov���Հ����݀����݋�ȱ�܋˔X�\�o����"�1�!�������텿����B��$|7��b�4����^�3��X�kp9��.s!xҲR��;%qLEB�4��gj��헍65
�ozG��._'�U�S�?q�:�m�B�83��zv�|i�Z��G��f{�;N����P�;���I@u4�(�E�o����5C�ǃ1����g�:�e j��R�H�k�J��'�5�$��r�=C.Y�'�e�<���r��%C(	��H�c�$�	j�Ӊ�~���&�)�YdI�%�Ӻ��|�T)-n,���,�%�G7�v�Ԥ�Ǡ����/]�86�R�� \~S�x5�[57���v��p;O8�x�;-s�4Y�r�fK�P��"�+!E�VB�}�O�+z}q[�T��N��~@C�?y���}?y�hl��Cd��(~� 8�	ƈH��[��xݱo����;^gk��wᝮ�3�߆v����~-��E��H�����"�_$[K�i|�m/����0}�f����>�3ۆ`�p�n���0}�f����>�3ۆ`�p�n���0}�f����>�3ۆ`�p�nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r�o�K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/�W����}�^�+���x>ܯە��r�nI���4��&��$���^ܓKےi{rM/nI���4��&��$���^ܓKےi{rM/n��r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�_*�ʅR�T��U.*K��R�T��?(���Z�nР��(?$���E7x0���s��ø��-���$G��Rߖ��]��d��w��%K~#�����0����D~9(P~N��-\�嫞ܵsۖ�{r��nZ���W=�j�-\�嫞ܵsۖ�{r��nZ���W=��ϊQ�iG.zR�_�K�mwc���$�)��T/��
���w�{�8��B�B��C;XT�s���qw�6��r�;���(�a�v=�Mɬ�m7�j笗�i�?�^��ߋ2_����+�+�,h\o�*\d�ư��X=�#������y_�M$�WЪV(<m���ɵ��q�b4�2�&S��Щq�\e��d�FY*Q�J�d�R����2�J&W�D���bڗض��-��J����R�$Լ�5/2����)�@Ю}hW>�+�Zϭ
�օs�B���\��w?2��̧s�)���w?2��̧s�)���w?2��̧s�B��С�6Hw[$;���I���nwM��I��I7;�&�q$���0��L?���+�����2�?�~���s�߹��nd���&��W���� ��(��J'�R��� ��.�J'�R��Ԣa�<d3��jQ��_��!���3R��jV1l�@R�������K:.4���K:.4���K:.4���K:.4�,���gkax��_x��cy'��<X�I���O7��,����,��Ě�h�YŏvX�`E�v�`����J�/�UR���@_Ԫ��P�*���T�J�/�Ua��i@XcJ�PҀ�Ɣ�4�,1�a�(i@XcJ�PҀ�Ɣ�4�,1�a�/���~�<o�G����/��/Ҁ��X�Հ�Ƽ�5�,1�a�xk�Xc^�C�
ܨP��B�7<hc�Ɔ8�ovߍ�ۋ��X�7��1��~�|hc��� /��,W����E��>�b�K�`.sX��oƕ����P9��iY)@Y����"�gi�3����K���.�����;�����<�����iϊC�7�� dlӷC�@䵵���\T7+��Y�l,�= \I���Ӿ�3�pj���Pzqd�#��@ꡄ��Y���*r��',��r� j�������r�<��Y '�5 k�z��@O>�C.Y4�T2��N4���P` T1�g��~��Mi����Ipt��,�
KA��=,���@K$�y��杸5(3���%��ǲ�P_�wH����n[5�e�o{x�l�6^6qʋ�;s�4Y�r�+��2?qY
,�E#�}q[��wE��i��b@C�G���_O�E���^@q����hn���i����D$! 7��o�-�vżn�gk��xa���3�߆v����~���;]������"�_$[K�i|�m/�-��E��H�����"�_$[K�i|�m/�-��E��Hf����>�3ۆ`�p�n���0}�f����>�3ۆ`�p�n���0}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r�nW����}��/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��N�/��K����;��I^�+���x>ܯە��r�nW����}�&��$���^ܓKےi{rM/nI���4��&��$���^ܓKےi{rM/nI���4���ʅ�r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�_*�ʅ�r�|\�_*K��R�T��U.*K��R��\�?.���v�1��z��qpa�/\;�Z�qG.{t(?�K��rD~94��?P^>K���ض��t��Fr��7=qM�j�(��R��nZ���W=�j�-\�嫞ܵsۖ�{r��nZ���W=�j�-\�嫞ܵsێ\��v�r�(�j�4����v#��R��-��{�� ܖ�8��{�rr�A�T+�%
��-|qz�8�w=���ޚ����e�G-�~#m��l�W�#��{Y��PYA\wtA�Y4�\o��\u���G��{Yds��H֕B��RLY$��M.O)��%}�l�Ƃ�xД.7��#���R�#��%.�#����hPx�N�)ԣ%z�L�R��Ԣ{��mK�[R�+ԡ%z�$�R���P�O��'���s�)���w?2��̧s�)���w?2��̧s�)���w?2��̧s�)���w?2��̧s�)���?�;��N��S���C�hP�>��)�@�2����)�@�2��̧s�)���w?2��̓��I���ne�)_�
W����8�^������Fw�#!��l3R���Fw�#;���J6�FŰzH�I��"ϺE�q�Z~�M )r�K�i�Y6���t\i���i�Y6���i�Y6���i�Y6���i�igEƖt\igEƖE��,�$з�"���-�H�o�E}�([�E�b�,Cqb��X7�Ɔ0b�1*�ī��dx߬���k��\g�߬����~�<o�G����Y7�#��d@_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�_֬�j�/�eB�vT/�eB�vT(cr�C�
ܨP���8�-q�W(��@_����P䀰�'����\>41�_�b�����#�^4��E��>�b�x%��4���\��J�o�+)�9��.s!xҲR��;%qLEB�4��gj����TmB���;�����<���K�J�3�]���A�7�= s���9����#�Ÿ������ ]��s�0�3�@�FD�f��,� uc�^Y�"4�5�>�M8C(	�d哖IUr�<��Y*����CP��jy\�T5P֜j�P��r�'�H	���5�ƜX��$@A�(��(�!�;����uA�4ဲ��E &�s�Ye<V�@�_��q�3��:u��ʹ��^�P�́xz�P6c������(��k"Ĭ�ř/��2^J�\�Y������]����ă ?T���i��cO�+��b?��"�~�/��"���hl��Ct��O�P$! 8�	ƈE�XT[��xݱo�-�vżnط���b�7[��x�0��~���;]�gk��wᝮ�3�߆v���_'~��ߥ�w�|��_'~��ߥ�w�|��nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r��W��J�~I^�+��%x?$�������W��J�~I^�+��%x?$������^�~��ߥ���{��^�~��ߥ���{��^�~��ߥ���{��^�~��ߥ���{�/~W������^��+���z^��Kߕ�{�L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��/����B��P�.T/����B��P�.T/����B��P�.T/����B��P�.T*�
��B�qP�\T/������D~.\e
�B��J?���nQ�䖮{}���-\��0~%/�Q��~9"��?�<|������1�R�x0��z�Њn���\}�9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>(�ϊQ�k�!��ʖ��K얩{��.�-T�寎&ց-|p���.J�B�o���O�~Q�nJ5+����\�5+����Om�Om6��%\�%\Gm��B֛��w���5��oj�!+��H���$���^��T�3���ixN�U�g:�OM$�%��䳿���w�0��ǿ���xԒ�Od�K,�idGk'��d�J]���a)��$�<l�����;�x��2��C0x�f߃������(I^�	+ԡ$���O��'�����I��$��~?�?䟏�O��'���s�)���p�IN��S��Jw?2�>S���nd���>S�����(|
�����~e?�O�S���� e?�N��S���~?�?䟏�M���+�Aw�Q=��O�3�������FC5(�f�ԣb�=$3R��jQ��J6-��E�zH�I )v2�c�~�Qb��;�>��"��.��"�;�8�����.��"��.��"��.��"��.��"�;�4Y�I���M}�([�B�t�,Cqb��ŜX�,��1g!�?���~� -q�R����~�<o�G��Ȁ��|�3�-q�P�~��3�-q�k��\g�Z�>���π��}B�5�q�P��z�\k�*�^�W�
�רUƽB�5�q�P��z�\k�*�^�W�
�רUƽB�5�q�P��z�\k�*�^�W�
�רUƽB�vT/�eB�vT/�eB�7*1�P��ʅnT)r�R>�P����\m�*�n�Wu��P�[��퀵�l�~@_��#�^4��x�>qX�X�����ج^�x��k
VS�iYM�e6�2�d/VJPGd�.)��Yƚ@��B�s�����*���U{�`ǣ�q��:�r�g�ҺM��M��C�H�T�e�x�Ф|�̎��Γ��,{4�?�,����31mC=8yl��C;rϧCP0*T5 j~Y�'��z��'�5P���T5�$����d�e j@֜iUjT5P�L	5�@DT0����;��,��Ӵ��w,w� ��ߍ��7�x�f{�:@�
G���A����_:IB�=:�Kpe\�yoG��(1��UaP�������@^e3�LX��س%�+���~.,��_E#�����ă ?T��i��b@{����b?��"�~�/��"���hl��Ct��O�P$! 8�	ƈE�XT[��xݱo�-�vżnط���b�7[��x�0��~���;]�gk��wᝮ�3�߆v���_'~��ߥ�w�|��_'~��ߥ�w�|��nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r��W��J�~I^�+��%x?$�������W��J�~I^�+��%x?$������^�~��ߥ���{��^�~��ߥ���{��^�~��ߥ���{��^�~��ߥ���{�/~W������^��+���z^��Kߕ�{�L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��/����B��P�.T/����B��P�.T/����B��P�.T/����B��P�.T*�
��B�qP�\T/������D~.R�;v#�r�T���K%/�I�D,����r9Rߔ~9%�H�K���ǻ80�����G*[��$�s����\}�Q����l����ϊ9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>(�ϊ9�(��e�^��r�Թ:p��T�9��p`��ϓ���-A��]��#���qJ5.)F�r�ԮX����znںo�x�V�_&;n�����s�Cslb���c���7�m���eH��_eJ�#�8�J���G���K$��M$�~��O����t[�7EƑE�i7�&�x�iOk,����O�'�v��Nֿ�����t��.�W��J��I^�I��!�]$3K���Q2�J&W�D�?RO��s�)���w?�O���$�AI?RO���$�AI?R���s�)��;��N�)���w8)N��S��Jw?���
���C�С�Ht%��I��$��~?�?䟏�O��&��I���nd���_�
W����8���g�3��+ԣ%z�g~߃�����.���C4�N�7���it��.�-��Ż[�kc�l|oԪ,C1gyg�q�Z~�M��d�E�q�Qgygw�qgygw�qgygw�qgygw�qg�"�<i-�Y���X�`E�vX�`E�vX�`E�v�`����`�_Ԫ��P�*�Y41�Z���Z�
�רUƽB�5�q�P��z�\k�*�^�W�
�רUƽB�5�
�ݐ*�v@����7d
�ݐ*�v@����7j벡~�*벡~�*벡~�*벡~�<j�_Ʈ5�j�Ʈ;<j�Ʈ;<j�Ʈ; -q�k�(\q@Z��P�‿���\�q�P����\m�*�n�~���Ʈ7�j�~�����|+Ƒ���@Y��>d|7��b�6+�X������*��xҲ�dt�s�
�2�+%(#�P�T,�M \v�p9�6Qbl�/K��/�P\~���mg�+�~�����W`���C������C�2^֟���<�����v�B�f$�H��)�@�n�Ā��` T7'N?I�@I�gP���	�$�1埖~Y��j��R�r��',�p�d�}8�q�gӃ j@��8�d���;��pH��mCl�wi׆@�H�H��|����W��v�������φ�_:I{⼱��
KS�G#T/P������k|ni�g�Ge��s��2^J�\��#�}q!tR>˧��\H2�N�a�Ā�[d�� !����#�~�/��"�~�/ 8��Ɔ�46@q����x����x�gk
�v��gk
�w��n��-�~E��ȷy��?"�wl[��v����~���;]�gk��wᝮ�3�߆v����~���;]�gk��wᝮ�3�ߕ��r�nW����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯے`��L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$���{�/~W������^��+���z^��Kߕ�{�/~W������^��+���z^��Kߕ�{�/~W������^��+���z^��Kߒ`��L�I��I0~I&�$��$�?$��A�(P~J���A�(P~J���A�(P~J���A�(P~J����rD~9"?��H��$G�#�����rD~9"?��H��$G�#����P�\T*�G����D~.Q��G����KW=�>��qJ?��bs�ܯ�����Qʖ�r�ø��Ij�Њn��ݞ�wz��qz��R��nQ��T��0~��9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>(�ϊ9s�\���>)k�9��(��e_'�Щrw!�>Ȥ+�l�W�YZ��G��p~�j����\�������Y){��=�9��q$U�!m�H<R�9C���ɚ��w�W;�/��K����S�
z.N��Qڹ��1L�_��E�?l�+4����W��)^��H՟E`E��Y�J��U�d]�4��Ɠw���gk'�x����kc��%z]$�K������S���pz�^a)ԣ%z�L�R��~ ����'�
S��Jw?�O�L��$�D�?RO�L��$�D�?2��
S��Jw8)N�)��;��s���pR��
S��Jw8*?�
���d�BY!ВM����I��$��~?�7?�M��s�+�AJ�R��&W����#;�����f�+ԣ;�x��7���it��.���E�[f�I��!�]$[���v�1n��@q�$�O!�[����-?k&��d���$.Y )rȳ���;�8����;�8����;�8����;�8[�����8[�����������������@_Ԫ��P���(�Հ��X�ըUƽB�5�q� R?��W�
�רUƽB�5�q�P��z�\k�*�_����[#�9l���?s����[#�9l���?r@����7d
�ݐ*�v@����7d
�ݐ*�v���#� ,�݀�?v���#�`,�݀�?v�P�‵��8�-q�k�(��@_��@�$�H�I���#�$
��*���#�`-q�P��#�^4��@Y��>d|6�b���ج^�x������*��@Y �Y �\�B��̅�J�J���18�H��\v,�h��k"Ǐ��U[\���|�C�ܥC�j֜��Zs�����3�s�7��H�W���Y��f�����ݧ>�;�!��"�K 4����-8�$T1Ӄo�H��1��=C8��ϧ@������@֜C.Y4�v�CZq�$�HӍ&���q$T1�;��N$��:��P�X�1�i_��%���� {�x��ŏ�3�@G$�0�!���R�b�i�r��0�w�=2AIj�H��j�2����@�x����v�8�x�;-%f",�y+��rZ|���Uą�H�.�\H:}q ��:-�+�m��l��#����Ⱦ�����ȼ��Cd 8��Ɔ�46-�D"�4B-�D!��*�¡��*-�~E��ȷy��?"���[���}ݱo�����;]�gk��wᝮ�3�߆v����~���;]�gk��wᝮ�3�߆v����~W����}�^�+���x>ܯە��r�nW����}�^�+���x>ܯە��r�nI��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��L�W������^��+���z^��Kߕ�{�/~W������^��+���z^��Kߕ�{�/~W������^��+���z^��Kߕ�{�/~I��I0~I&�$��$�?$��`��L���A�(P~J���A�(P~J���A�(P~J���A�(P~J�#�����rD~9"?��H��$G�#�����rD~9"?��H��$G㒅�r�T��?(���#�r��\�?(���Q���ø�M�j緧ⵊ��b��շ� �pa�.�Sw�ݎT��[_Ȍ�Q��T�嫞ܵs۔~9%�IG㓃�w����r����G.|Q˟r����G.|Q˟r����G.|Q˟r����G.|R��n9��i��׷�K��Է��[C�q�n#o�������^9~w�8��>H�.d�ܬ����nZ������!�G��mվ۫}c^�-�/n���G+�w�~[���kY���O��w����>P�G:�*v6I�RZ��x�T-�7d�v�YߩY����2��(����x�ȷ�,�w���O��+�]$�R��`���.�W��w�u�M.O)�dҞ�M)�dҼ�W��J�{	&$Ԭe:�d��I)ԣ$������jV2�J2S����Q�+�m
�d��Y!�H|e�d��Y!�H|e�d��Y!�H|e�d��Y!�H|e��$�AI?RO���$�AI?2O�L��)��;��s��nq�M�6W����)%�N�JǿR��`�����E�����_���=�[K��iu�m.�@md�k'�Y>�ƖE�i4[��E�Y��Y�5�������~�O�`t^��݃�{�b�1*�0Ī,��[�ȅ��[���Ī,C����~�<o�G��Ȁ��|�3�-q�P�~�B��U
G�H+� X���H��#� ,��X��B�wj+� R_r@���I}����%�$
K�H�ܐ)/� R_r@���I~)�v�ې,Wn@�]��v�ې,Wo��~N[%�9l���_���~N[%�9l����ʡb��ܨX��B�w*��T)r�R>�P�}˖�~N[%�9n+��q]�[����W�����帮�-�w�
K����)/��s�W-��[%��@\V!qX��bG�`,��ŉ�>d�~�x����%��9�@\�3�ߍ+)�9�����ҲR��;%�H��1�x��"�qܨ6R���G���.?�P}&��y��l��Pl��>Ȭ�q�3�a��)zv�Cfe|桹�r�P�="�ӿ�=Pf !��E�WӃ4X�g�5C�H�;��q`"��:Ӄ z'N&��t��@��'N$�t��OP�N=C\��H�N$�0 ��Dt��h	�T<	�
@�Y�I�='i�ON�d��>Ο�r�+��vI�iky�^����4�Q�e�N��wH��2~5@�ŏ��x�ر�l����YƳƑ�h�+1�9�ŌVJ���� !�@~���M�a��[V"�b� =����b? !�������Ⱦ����46@q����hl��Cd 8��Ɔ�46@o(y@�x����w��n��-�~E��ȷy��?;���gk��b�7l3������x?$�R���������/�K���������/�Kߕ�����W��J�~I^�+��%x?$��v�0�׆���;^gk��xa��3��`��L�I��I0~I&�$��$�?$���{�/~W������^��+���z^��K���x{�^�ׇ�����x{�^�ׇ����{�/~W������^��+���z^��Kߒv�2N׆I���;^'k�$�xd������{�/~S���t��N��)���:^��KߡA�(P~J���A�(P~J���T��-�%Kn�R۲T��-�%Kn�Rۈ�rD~9"?��H��$G�#����T��-���$G�9sێ\��=���n#�r��\�?(���#�r��\��IG�9R��E7c�2���Q���8��or��(������C������?��-��j]��l�䖡���?�Z��KP�Ij�-C�%���N)�އvpn{�������J5+��k�B�p�6���>ܣR�K_R�J����`�2��o����p�`�p��H2��m��k�"�}
VIPmJ#����q{�:���rr��ܞ��/�{^!��`��_=ҜJv�Yӵ�������|W�����_(\��Wq�v����:�Sg���ԩ)���+_�6�d�#�\����K�w���С�p���X:�E}�(��B�t���W��&����k	����Yd�ƑP��*���������W����{	&�a$Ԭe?�O�I�XI5+&�a$Ԭe?�O⒅s��\�hW8��6�s��\�hW8��6�s��\�hW8��6�s��\�hW8��6�s��\�d���'�
I���~"d���'�&I���~"e;��s��nq�M�6W����)%�N�JǿR��Ԭa�=�3��`�m.�-��Ŵ����_����]|�����O 6�}?�,���h�k"�v�)Ƴ�k=?y���04�������=���`ŘbUa�TY�%P���Yb�E�bU=��7�#Ɔ4�o�D�j�Z�>��`-q�P��z�#��
G�H+� R?�@�d���G�T,Wv�b��ݐ)/� R_r@���I}����%�$
K�H�ܐ)/� R_r@���b�r���+� X�܁b�r���+� X��-����K�r�/��d�'-����K�r�/��d�$�I~)��R%��
K�H+� X�܁b�r����/��d�'-�w�n+��q]�[����W���"K��/� R_�@��-�a\�9�t���3�B��
�%�
K�*��T,V/P�X�����lV/d�~�x�������`.sX���cƕ��VS`.s!T)Y��d�dvKƑ�X�b .)��EB�Pl����{�<�A��z���5+dm9�ҹc�o�.�@��n�ā�G�,�%�&�qM8am@ӆ�r�'T��It���(�@���@����5C�Dt��i�3�@E�5P�@��8�'�1��Ӿ��F��t���P���0f !Ӊ {N�����P %�iڅ�wIt4���0V����b���@G$�yqԁ��/N�p����9c�Sӯ�P���-��
e�hY��}�X㵱c��x��*⚟Ge�Ĭ�B��+d~JⲄ��Sd� ?Tض�Ű�b-�+�m��l��#����Ⱦ�����ȼ��Cd 8��Ɔ�46@q����hl��Cd� 7����x��y��?"���[���w��n����żnط�� 7��o�����{���K���������/�K���������/~W��J�~I^�+��%x?$����������;^gk��xa��3��v�0�׆I��I0~I&�$��$�?$��`��L�W������^��+���z^��Kߕ�{�/�����x{�^�ׇ�����x{�^�׆W������^��+���z^��Kߕ�{�/~I���;^'k�$�xd�����v�2N׆S���t��N��)���:^��Kߔ�{�/~��A�(P~J���A�(P~J��R۲T��-�%Kn�R۲T��-�%Kn#�����rD~9"?��H��$G��R߲T��?��H��n9sێ\��=��ϊ9s�\���>(�ϊ9s▮{r��o� ���5�4*\+� �J5.��Ѐ\�4>�$�ܲA�(T�Wz)�B�º��;o���ö�0�;o���ö�0��s�sܔ~985+�r�\�%��ܵ��E7zp��\;����-\��5+��������o��Ї��aݞ�'���,�����r�(R�J��6��R�)��([Ȅr��p�6���$sy@����3�J�|�_=X�V�U�UoUX�S���Y�5��_X׾?��{W%�n��<.W#c����p�NRb�5�VE���8��X�!\���E��k�Y���v�.��"��ŝB���Kʺ.5~��������M$�T-�k�)�d�<�I���<�S���u)=
�aB���T�%:��S��о+�U+%����cd��Y>,b7:H�Β#s����"7:H�Β#s����"7:H�Β#s����"7:H�Β#s���Fо"h_4/���6�s��\�hW8��6�s��\�(W:IO��S���jVMJ�I�Xw�,!��|3R��jU�lO���lO )rȶ'��d���$.Y��d�~�M��d�~�M 8�rk� 6�:U��]�#��dt[̎�y�}��gݟ}��҅�Ɣ-�4�l1�a�([iB�cV,~�b��^,~�|j�Ʈ5�j�Ʈ5�,�݀�?���څ���,Wr�b��ܨX��I~)��R%��nsr��˖�7.[�ܹnsr��˖�7.[�ܹnsr��˖�7.[%�9l���_���~N[%�9l���_���~N������g;�#9����H�w�Fs��3���%�*��R_��I~J�%�*��X��B�w�
K����)/� R_�@���I����%�$
K�H����+��0�[�ºD��Hs@�,�P���IzB�b���ج_��b�6+�X����%��K��sm���b�J�w�+)�4���\�B�R��J�J�엍#���@\S�g���<o�P�]�-�ڂ�*�����j
V��s��rǲߧ>��QI:w8x4�YhR>�~V@M 8�3P�H�*�N�����>;�M��N�b���2���5C��Ӻ@�8�w��:�1D���q��@G uc�]8�'��N<��2�� ~��G�0ӵ������P}�Y�G��X�`�tP��~Gr�B��v�Cw�Zu�T����,ziU%�R�����E���x�ر�kanq��T�51bVgans��2^J����d~.@~���M��l[V��b�����u�@C�G���_O�E���^@q����hl��Cd 8��Ɔ�46@q����hl[ƈE�h�[ƈE�h�[���w��n��-�~C<nطy��?"���[���xݽ���Kߕ�{�/~W������^��+���z^��Kߒ`��L�I��I0~I&�$��$�?$���{�/~W������^��+���z^��Kߒj\2MK�I�p�5.&��$Ըd���R������W����~�^�+��ex?l�������W����~�^�+��ex?l�������W����~�^�+��ex?l���}��/�S���t��N��)��e:_l�K��}��/�S���t��N��)��e:_l�K���b0~��#���b0~��#�T��-��K~9RߎT��-��K~9Rߖ�{r��nZ���W=�j�-\�嫞ܵsێT��-�G�Q�䖮{r��nZ���W=�F�(��%~�����\}˃�pa�.�{s�C�����4�W�-|p� ��8�΃��¸7=��~Z������X�΃�Ѐ\��Br�@.]ˡ �t .��ӊqw�6寎j��-|p�`��\*��G ���7�k��!Q�?��އm��Q�<+�߈��%8b�[}��~�J�V,����{���5��l��Q_�����b��'K��]�_��?��%HnB۞��+��zۤ�硹���W�4��E�V�U7�)\��K�-������[�.��:���K�����[��tR?n@{�"��O�`E�c��WE��t[�4��H��i4�ƑP��-�k�)���z\�I��$�<�I��%:��S�I�:��S�I�:��S�I�_�/��%���s��\�"0��Β#s����"7:H�Β#s����"7:H�Β#s����"7:H�Β#s����%?�IN�)�RJ���$��I)�RJ��Ō��c)�X�5+	&�a$Ԭ%x=|���jU��J��WŰy<[�Űy<���$.Y )r�K�i�Y6���i�Y7EƑt\iEƳ��ҭ?�*��Ү�y��o2:-�DY�gşv|Y�gşv|-�4�l1�a�(��Ջ�X��Ջ�x��׋������쀲?v���#�`,�ݨX��B�w$
K�H��)/� R_�@���I~.[�ܹnsr��ˤJ;�+6�D�ۃ)�R;��w$H�H2�ܐe#� �GrA���)Y�R���gJ�2��0e+8`�Vp����)Y�R���gJ�2��0e+8`�Vp����,�~@����w�9ߐ,�~@�����2%�yns��s��[�¹ns
��+��0�[�¹ns
��+��0�[�ºD��t�Y�)@岲�ed6@��l�g0�������%��K��,���Y/m��^?P��mB�m�9��)YN�R���J�o�+)�9�����ҲR��;%�H��1�x��"�:ȱ�k ,,�r�g^���mA�x����:u\��c�!��/SӞ峤�8t��ꖝ���,��+/8�o������<���uA��Oӟ�ޝ����� ���*��p`�T(	p��I�P�@��T3�=�U�f�=8�p�چpE��!���:O�.�����?pf�/Gk���E��r�+ r9����K�.�>��vʃ�Wj�!�?�;�9zd�A���}����Ŏ;[x���r��q��vZ��D-�r�+��2?�W��Sd� ?Tض�Ű�b-�+�m��l��#����Ⱦ�����ȼ��Cd 8��Ɔ�46@q����hl��Cd 8�ط��x����x��y��?"���[���w��n��@{�R�
��T[����x{�^^��+���z^��Kߕ�{�/~W������&�$��$�?$��`��L�I��I0~I^��+���z^��Kߕ�{�/~W������&��$Ըd���R�j\2MK�I�p�5.^�+��ex?l�������W����~�^�+��ex?l�������W����~�^�+��ex?l�������W����~�N��)��e:_l�K��}��/�S���t�����A�hP~���A�hP~��#���b0~��#���b0~�K~9RߎT��-��K~9RߎT��-�j�-\�嫞ܵsۖ�{r��nZ���W=��K~9Rߔ~9%�Ij�-\�嫞ܵsۖ��R�;vZ�n�P��\;����ø�p�)j�ފqw��|��z��nxcې�w�ۖ�8z��=��nt�\��N)�Ѐ\��Br�@.]ˡ �t .��Ӈ\���_��z��Ӈ\�0.�:�޹�Dx��!�¥_���Ըx5.]χ��G �ض��������\e�]�T�B�Ix�+�R��5�~�o��2m>GShPŷ�Ə���GS���R˼Rk�$W�ȝ��
���#�nB��硹����4)��mH;wm��ƪA�J�e{���;�wY��q9W&����%�E��׾r��ߑl����b�>G�J�YT��i��=?�g 7�(gy"�x�+&�Md���)vrN�W�����9^�g$��RLE$��R�JM$��R�JM)ԤҝJMB��P�%�/�e��ad��Y.vK����ad��Y.vK����ad��Y.vK����ad��Y.vK�����S����)%?�IO�S����,e?�O��I�XI5+	'�I����Ry^�'����<�W�I�z����w���f�&�irhf�&�irh�k"�v�(�k"�k9Ƴ���~�O�`i�iWE��跙��>,���ϻJ,���l1�a�X[j��cV,~����_Ʈ;<j�Ʈ;<j�Ʈ; ,�݀�?v��څ��T,Wr�b��%��
K�H��)/��s��-�n]"Vm�Y��d�'H�w�Fs��3��2��0e+8`�Vp���)�PR;���wmAH�ڂ�ݵ#�j
Gv���)Y�PR��g�AJ�ʂ���+?*
V~T���)Y�PR��g�AJ�ʂ���+?*
V~T�����J�Α+?:D�����J�Α+?:D����!�%dC�JȇH�����:Fs@���g4�+""VD:D��A���r�Y岲�$t_�H�-��~[+"�9��,��P���B�k9�T,�P��mB�m�9����T)YN�R��dt�dt�s�
�J�_�+%(#�^4���\SqLG��b<n;x췍��
�lzE@����.?Q\~N��kN��W,x��u�t�ӟ>@�N��,�L���@p0f��@ӆ�r�yo�N�����.��x54�(���9B��NC}�	��
��l
��lZ��(	��9e���t�9�~��:OӯT����\��0��@M�f{��,�t��j�n�Ϥ�1������-��s�)[$t�>F��Q<DY�w����Şc1Md-�2�bVgbĬ�E�VJ�2?�WE\HR�M��l��Sb�b�����Hu�@{����b?��"�~�/��"���hl��Ca�4^�E�4^�E��6�Ca��6�C{�ȇy��"��C���w����!��D"���[����T��B���?;�^�׆W������^��+���z^��Kߕ�{�/~I��I0~I&�$��$�?$��`��L�W������^��+���z^��Kߕ�{�/~��A�hP~���A�hP~�S���t��N��)��e:_l�K��}��/�S���t��N��)��e:_l�K��}��/�S���t��N��)��e:_l�K��}��/�S���t��N��)��e:_l�K��}��/���A�hP~���A�hP~�#���b0~��#���b0~��9RߎT��-��K~9RߎT��-��K~Z��KP�Ij�-C�%�$�䖡���?�9����n{��~Z��KP�Ij�-\��w���ø�p�/\;����ø�p�)F��އm�c۝˽�훐{�Z�~K_=8���-|p�n{���n���}ˡ �t .��Ѐ\��Br�@.]w'N�й��aܟ8����ܶn|��^w$ ��Ǹ�q�(����v�'���Yb>�W�V;��7�ƧW�}l7�^D�o���b^����[e|�?�����e�׼��?R���[b��,^�Od��)5�ri�Y�p�C@�(�T�d"�g��"�J�����n���}7��oV�bT�ٱz�d�*9�K�nD�����Uɖ�R��ǣ�sCܡb����Sanq���-�w:/�D-�%Qg���Co�Ͽ�����r������p;�\��W�����9&"�`�)&"�`�)N�&��RiN�&�|K(_�Ĳ�s��\�,�;%���s��\�,�;%���s��\�,�;%���s��\�,�;%��I�XI5+&�c$Ԭd����R��jVMJ�I�XJ�z�^�'��R~�Y߃�;�yg~,����<���C4�43K�C4�4[��E�Y��Y�5���Y���?y���0:/vE��跙��>,���ϻJ���Յ�Ƭ-�5b��^,~����_Ʈ;<j�Ʈ; ,�݀�?v���#�j+�P�]ʅ��H��)/� R_���7.[�ܹnsr��o�J;�+6��GrA���)Y�R���gJ���ݵ#�j��<S��Oʃ�?*��<S��Oʃ�?*��<S��t*��t*��t*��t*��t*��t*��t*��t*��H�C�
��"�D*�T>)�|R!P��B�t*�t*�t*�t*�t*�t*�t*�t*��HmAb�ڂ�!��Cj
GE�
GE�
GE�
GE��GP �GP �GP �GP:D����:/X��H��H��������������������ꅜ�jsm�)YX�)YX�R�� R:�dt�dt�s�
�J�_�+%(#�^4���\SqLG��b /�����K��[PPc�^_�x8����EC���u��</Ө^��^����\����Zs��T7�x�f��@Ӈ���Hs�uA���Ӟ�I�%��~��e�3�r�Rr�U$�4�ӴF��1;��-t�P�����(7N����j�?��3��`#�{�J4��w��g��4��A�?ew�~�ܶKI���H���.^��ދ��Şc8�-�2�fGgbĬ�B��+qYB,��^������,��Sd� ?Tض�Ű�b-�+�m��l��#����Ⱦ�����ȼ��Cd 8��g��x�xg��x�xgy�w��gy�w����!��D;�ȇy��"��C���w��g���?"���[���w��������{�/~W������^��+���z^��Kߕ�{�L�I��I0~I&�$��$�?$��`��L�I��I0~I&�$��$�?$��`��(?
�B��Р�4(?
�B��Р�2�/�S���t��N��)��e:_l�K��}�(?
�B��Р�4(?
�B��Р�2�/�S���t��N��)��e:_l�K��}�(?
�B��Р�4(?
�B��Р�4(?
�B��Р�4(?
�B��Р�1?F����`�1?F����`�1ʖ�r���o�*[�ʖ�r���o�*[��~Q���7=�F�(������sߔn{�ώ���sߔn{��?�Z��KP�Ij�(��R�>���ܸ0��r���\}˃�pn{���n����\C� ۀ��T-�_���@.R����J5.�&�!�7`;f�Br�@.]ˡ �t .��Ѐ\�p��=��rw�;x0xT�K�J;Z
���>�d�G�;ȼ���p`�-R��46Q�V;�l\C�J�~�CkN�|}�/s����YK�2�*������p�[&s Ş�+(��_�y(xd~Z=���n�=�u��_>�d�%��O�E~���'����o�;p�3���+!
�pɑ4^T��ڳ�jη�}o^�v��z����k���n����hT�KI��*:m�^���H�q�)Nۀ�;�,I~(��T,�V�}/ϋ2?#��%]�"�`�<l�������p%z]��K���vrLE$��RLE)ԤҝJM)Ԥ�/�e�Yd��Y.vK����ad��Y.vK����ad��Y.vK����ad��Y.vK����aB�XP�V*��
�aB�XP�V/���|�R��u)<�R��0yd��J��9^�g+����yg~,����.M���n�E�dQn�E 8�r�g��04��E����=���`şv�Y�iE�v�-�5al1�a�X��׋�x��׋�����#�`,�݀�?v���Gܼir�����v�.+�P��%B���
K�Hs� Y���g;�����Y��egH�ݽ"Gv����)�PR;���wmA⟕�~T)�P��*��UC����!U�B�8�T>q
�|�P��*��H�C�
��"�D*�T>)�|R!P��B��H�C�
��"�D*�T>)�|R!P��B��A�
��(�P*8�Tq@�<�/Py�^��HmAb�ڂ��z���z���z���z���z���x2��2��
��!��CzD����)�,R�X���H��H��������������������ꅜ�d
VV$
VV$
VV$
GV�
GV�,��j)e��̅P�f/ƕ����/Ge`.)����#��16q����:���\��k`���A����&��zeA�1ڇ�e���[��A�>�{��u.���`!�k�;Y$�r�),��j�x3P�i�P�x="���P^�����~�|�O�(N�3�t�?���9��A�,xdTsN[�5k�3Qc��?|	���3+�0пP�x���:MӊA��r�Χ^)��1څ��*�Y�Pc/ag�,�;�?8��Y����[�e�̎�ŉY��2^J�����WY�Yz(bA��l��Sd�����E��b@{���m��~@C�?y���}?y�hl��Cd���/���/�!����!�����P;�jy��"��C���w����!ߥ�C;XT3��E�h�3��w����I�p��~�^�+��ex?l�������W���5.&��$Ըd���R�j\2MK�I�p�5.&��$Ըd���R�j\2MK�I�pР�4(?
�B��Р�4(?
�B���t��N��)��e:_l�K��}��/�S��Р�4(?
�B��Р�4(?
�B���t��N��)��e:_l�K��}��/�S��Р�4(?
�B��Р�4(?
�B���*[�J�����d�o�*[�J�����d�o�`�1?F����`�1?F����*[�ʖ�r���o�*[�ʖ�r���o�j]��lF���v�j]��lF���v�>8c�2��~Q���P�Ij�-C�%�$�sۖ�{r��nZ���W=�j�-C�%�'����t�R�K��Ɔ��=_�_��z��k������,��RyOy�����^�;o���C�����;o���C����;������>���S���)[-��k~�B�����ub���Ы�m��[�w�ޝ.�%�Q��dW���ȸ��6=��g���f�}CdHc)��$>�m<�ݦ��\���?%�~W��e�^�{�v�|Rk�R+�)�)�Ri�H�r'%��D�;p��}���Ფ*��f�J���6]�t�_Jv�{��z��ʶ��z��K7*/��Oc����J�)�wdY��x[#�bVv��Y�s�N�K�����O��R��U�eP��Uߥ���x=�^�����MJ�I�Ȥ�<�S�I�:��S�I�_�/��%���s��\�#�9<r�'�\��˜�9s��.rx��Od��Y.v�Ō��c)�X�4/���J�#R��|Wо+�_�/���|�R��u)<��I0yd�K�J��43��irn�Y߃�!�\��ɡ�\�-�Ȣݬ�-�ȴ�������Ү�y��o2:-�DY�gşv|Y�iE�v�-�5al1�a�X��׋�x���������#�`,�݀�?v�b��6+�q]����\Wn�u
K�T)/� Y���g;����s��eg-��<�Vp���$woH�ݽ"Gv���$wlb��e�~Tq
�,�PY�*��H�Ag���"�D*�T)�,R!PX�B��t6��t6��t6��H�C�
��"�D*�i�q@�<�Py���A�
��(�P*8�Tq@�.�Py�^�
A�2�(�E�8��q�<�/Px�~��H�A�����ڃ��ڃ�#��VCzF)��7�b��2�#��8���)m�,��$t�H���H���H���J�āJ�āJ�āJ�āJ�āJ�āJ��B�Չ�չ�պ��Yj)e����P�f/ƕ��#�^6)%@\�+qLD�1�8�E�Mxd�x�.[P5�e;�e��j��T/#T<��TJ�?���U>X������ޥ���� ds� nS�����Xg�3��0f��@嚡x<�rޏN�%� ��v�x���gI�u P~)��=^�8ymsj,tuşn��T7�0fe|�Z����Kӷz�oz��,{�eҺD���#H�������GE�kb�����*���#��fGgb�s��2^J��~/��$-?�e�ă ?T�����6-�+ql1X�a�Ā�[d�� !����#�o�/���~�/�!���w��g��x�xg��x�xgy�w��gy�w������P;�ȇy��"��C���w��	^�ߥ�C;XT3��w����I�p���W����~�^�+��ex?l�����(?
�B��Р�4(?
�B��Р�4(?
�$ԸhP~&��$Ըd���R�A�hP~���A�hP~����}��/�S���t��N��)��e:_l�K���b0~��#���b0~��#��}��/�S���t��N��)��e:_l�K�T�hP~�#���b0~��#�|p�>8l�6O�'�s�9���o�`�1?F����`�1?F���� �q�>�r���o�>8c�2��l���(��b0~�K�#�����Իe��R����\�+�s�����w=�j���G.{q�IF�r�~98?������s����}��B����=px�Y����6}P��A��+I*�R���P��UJZ�������~�N�Ӈ������'z���V :�~KTy$��΃���D=��=���J�D����>w8l����8�K����[�F[�!J�]%>J����	K#J��M����.2߳ȹ��a�f�+��S/�n�j�$�
ƾ{vN�qW���U�*�z�'��X�K)b�,\����r�8dN���f��~Y�,�6o�R���N?�V۫/N�[�� �a��U�p��p߲�l������E�W/c��u�{~��$W�
}|��8,[rE��'Emżm�&�)Բ$�>k� 8ڲ�ĊS����yd3��J1tL���\�=qJN�z7�����R�J#�pa�)G�M(�I��)4���iu��c )v2k'�T��ʔ�9R�Y>$VJ���R�Y*Rk%JM)Ԥ�LE߃�;�yd3K�C;Yd��ɢݬ�-�Ȼ�\���`�<l�y*�w���y*�x�0�-�dH�~������]1��C��K��it_�(�\j���1^ȱ#�|lWs��w<lWr�~(%��.+�P��%B���
K�T,Wƒ��9္�B���
Vv�)Y�P�gl�H���ߒ#�9n)
帤+�␮��D:Fq��C�g��D:Fq�.�\��mAp0�2�"�e�P �8���q�,�/Y�^���g}:�+u�V4뀬i�mӮ�P|�N��A��z��!U��*���?��?P\7�b����	��J�?� Y��p�9�i�+u��`�8��qm�,��PY�b����Ag���+u�V�����xo-�-��������xoH�-�#�����8�H�#�#����.?P\�p�[�[d�H)N�,R� R:�dun��������/�#�/Vb�,�� ,�� ,��E�����",�h[��|o� ].ϖ�o-���6����'PR�F�)-ZӨ6���IB�>X���c�sӞ�.@�ky
��9+�x�Yf-� �Ź��gǐ?zX3~7�j��3u��7P�3u��5`Ɯ0A��8am@�?�q�E���L��9d�$G7�&�\�!����E ���Ǌ�P��䵺�mk�ty>���*�텾>�,�?8�tR;S�b�i+4�~s��^J��\���qr����Ֆ�$����6-�+ql1[�}��g�m�}��g�m�}��g�m�a��3G��t_���;�l3��ž�3���;�l3���������P%}�C�Ơw����+�b��!+�bM.$��R��!+�b��!+�bM.$��RM.)��%8?��������S��Jp�N�)��"5.�F��(Իe�lF���v�`�1?r���o�*[�ʖ����d�m�*[vJ��
�B�vЪ]�*�m
��B�vЪ]�*�m
��B�vЪ]�*�m
��B�vЪ]��l�Rߖ�[��K~Z�o�U-�j��-T�媖�F���v�j]��lF���v�j]��lG��#R�Իe�l�Kᖩ|2�K�Q�v�.}�˜*��P�t��B9R�G ���#s߲|p�>8c�2�K�Q���0~&�~��ߡR��?*�󿼏�?�{��R�|���9���}f�
��;h\ko��������m����>�繧�(�ϒ,����,g3�Ӻ:T�KE{"5�6Q�)޽�C���)��Z�H0��$�&k5��*��R�(\ƠT�=��I�H�)_���5d���w��m��X�d>/�p���C`���;�=M����`6���]7c��Yd�E%�r�-�x�Ǌes��PIg7zJ�Xd�~��4�	g���K���>��e�����ߑQ���ȍ�e��%��O;��w)<�Ryܤ�I�r���'��O;��w)<�Ryܤ�I�r���'�$��I��nK7��"pȜ2'n�t	U�܋��*��YzƽZ��Y�^P�]����\��y'�ߞ�~|�������ܼA��e��Gpzp���/s�oŵ�o~�w�*�rI��KP�W�)&���ȍ�MB��,�z�_y"�2?",��|1*��v|�C���v>�t�#�J7;8�JEd�I�:��W��Ŵ����_ߥ��)4s�9��H��+'Ċ��"�T��LE$��]�<��ɤ.Y )r�?k&�x�h������C<lg���%Qn�U�%Qn�U�"�6D[�Ȑ��?y��{�:/wdY�k�PƯE�ҋ5Ƭ-���c��g���xخ���PK�@Y/�P���B���
K�Hs� Y���x`.s�P�gmB���
Vv����)� R;�␮[�B�n)
帤+�g��D:Fq�.� Y�C��[�P9o@�7�p0ޑ�G�ˁ��?�8�H�#�#�����8oH�-�#����[���o�8uC�4���V*Ǐ��?P�-cN�:��Z�A���2�m��8��ρ!t��P�t6��C��mAqՎ[�E�nq�>�P|b��
uA���)��St��j8��� \:@�āp5����:GX�c�p5���[zG��p���#��G����� X��@�Jt�b���)�GV�,���Y �Y �Y �,R��H�Ƒ��҄�҄�҇��IP�8�E�-xO���,��ځ��/��`ǣ��9~��� ˗��=sL��v�)�w�=�=:���iϮ� d��ӴG� nI�dJ�_�^�sf-�*��4Y��&�><�gǀ�,��E�@�E�@M��2�qP�3#�%�d�����N���N޸<=8|����8�IB�9�����T<���/Z�.?'�|��([��b����gE�e�,S-�8��9�H	/%E��J@b��f���5ŗ���d� ?Tض�Ű�n�[a�u��[a�u��[a�u��#��1�����t^W�Ce}�6-�E��6�Ca��7�Ơw����+�b�5�Ơw��	_k���	_k�ip�&�
���	_k���	&�
�ip�&�
������S��Jp�N�)��%8?������H?�R햠����Z���5.�F��(��e?r���o�*[�ʖ�r����*[vJ�������d��|p�>8l�6O�'�
��B�vЪ]�*�m
��B�vЪ]��l�R����媖��Rߖ�[��K~Z�o�U-��K�#R�Իb5.�K�#R�|~D~?,�>��϶9��-T��0}��ߖ�8c�>���d��,���r��p�F��(Իb7=�'�s�9��(Իe�l��mw�X�/nW�!T-�����]�*ɼ�@p��+�R����F����ގ߻���:�m+jK�#%9/X��U��B���ϗ��I�l�-?"�)K��_)�n����K����Ξ�+K�j���OEbǥ�JY�V����V,ؚv�>��~�|�N^;,��d�+c�xc�l�XV������׼������;�M�rX8��m��j;	B��JZ���u-_l�K.y{���)p������'B��'ͫ,�a�p���,�8�ۆ$�E��g�Ȣn�I�$�2�?e�щ���,\����r�.R��X�K)b�,\����r�.R��X�K)c�E$��K7%����f�8dM����f�`΁*��v/�|J�^�cv�;��7vr�.$���m��-gkY���%�Z�YmC��\�M���}�~.����������w=ߜ;V#rP�\��+��;�O볃R�z�$�-���������Y�e�����_d��P�%�J���R�Y>$Qʔ�9R�G*R(�JE�H�0{:J΅R��T�䚕���I0y��w�R(f�&�irhf�&���-?k"���h��&�\g���b��-�dH�|��g��|[�Ȑ����������,��f݅��dY�k���k�ȱ#�|lWs��w ,�′_��I~J�%�*��,�~@���[+8yns��s���ߒ#�$
G~H��帤+�␮[�B�Fq��C�g��D ˀ�A�@�.P\6��oH�a�#���\t^�mAqՊ���V*��TX�.:�P\u:���uAq�����S�灦��eӞ˧<7N��ޝx��:���u�ӪV�륦��@�t����ρe劁e�xYM�A�.��s��H�)���:u��0e��:Gm�.:�P�:��uC�4��i�������? �? ���8
wH�)�#��t���8
tp�2�)�e�S�ˁ�A�X�.�\b��p5�2�)ܷ8�����s��-�+u��,R�P�K-B�,�4���i!x�:B���.��B��B�b����I^6q����:���@_i ].ΡT�x��[���GG��)[#i�sOӘ6ݧ>)n����2��`���;N{�KT��G8��!�;DR�ā����I�������:>�����#�#���	e|�9&K��)���2�����It�}%à��t��=}G�<U�:��u+c���e��9l�T/��t����kz.� 1MOE�e����s�D[��$����W%��
�,��ԃ��H2�M��l[V��b����Ϻ����Ϻ����Ϻ���f����~��/+�!���������!�����P;�j�@�������P;�j���J�X����I4�T�K�J�X����J�X��K�I4�T��������S��Jp�N�)��%8?������H?���-|p�_2�����-|p�>8c�1ʖ�r���o�*[�ʖ�r��d�o�*[�ώ��s�9����|p�>8c�1ώ��s�9����|p�>8c�2��'�Q���7=�F�(������s߲\�l�>�%϶�s��}�K�l��Y!�N��d���>8c�-��K~Z���P}��K~#R�\�e;�m������7=�]�o�s۔a�1˟lr�����5.�F��-R�e�l�K䖪[�������v��N�@����_�#��+��m�{�.�.��v�;��:��S�:�_/1�VA�qL\F��c�Y}Ď�ʽ\i*����\�(���/������6�?e��d�-��-+�#��B�����%rc���S2�0đ�l0d�&M��q��>J��t���zݚ�M�����KL�edY���:Û2���� ��m�2����Onl�K������Y�t�Q:�
N��k�&��dN����h+��T�Rhʶh���|Yܥ���r�.R��X�K)b�,\����r�.R��X�K)b�,rH��_�f�rY�,�2'��&rI��'���`�!��J���3��U�G�T�u;� �$�rd���ĥ���v΀��T�Eخ����+��]����H~��q����p|5.N�����;��l���w���&�a�e�1�X1oM)�X����&"�T��,j�*�\�;�<��"#R��T��U+:J�I�Y�0y�R��`�)^�g+����\��-��H���Y�5�[��E��T[��HvD��g��~������Z�KO�ii��~���a��[�܅��ȱ\qE��$~�xخ���U9�H�ې)Y��eg-��<�Vp��Y��$woH���"V~A���r�R�3��H�"#8�A�@�.�\��mAp0ڂ�a���j����?P�<~��x�Ax���������[jǧT�N�xY[�xY[�?�P~=:��z�A������u���ǭ�M�:B�.:B�.:B�.:B�A���=7�!eoN�Y�*��˧>��>��5�5�],�P\u����.�t����Ix�A������zs�H\���ycǦ�ǏM���<��<��t��t�P|u6���mA��ڂ㩵�Sj���M�>:�P\n���ApApApApApp2-�+|�8�����s��B�)���,R�P�K/�#�/GHP��\Sdt�P�IJ�b����J^6q����:���k<n;eP�f������j��(1��/Q\�f��l��U�>��vꃃiPe��/A�>�z��0�3�> ������A����4���4��Ӵr�7d�$�$|6I n�#��$~��?�;DP�!�%��Iw�zs����)�_;f�B�:�Tyc�]�?܇PR�;�::�H�r�����*�����|}��lt��Y 1MN�#��|��Ź�"��X��C2>R�d|��^��A��l��Sd������>�t3�C>�l3��>�l3��0�~�#��t_�����l���ž�3���;�l3���������P%}�C�Ơw����+�b��!+�bM.$��R��!$��RM.$��R��S��Jp�N�B�vЪ]�*�m
��B�vЪ]�*�lF���ᖾ8e��k�Z�ᖾ8c�1ώG�Q��~9%�IG�Q���rD~9%���sߔn{��~Q���7=�F�(������sߔn{��~Q���7=�F�(���$�sۖ����?�9�C�#��H�?�#���hP�?���C�hP��;��C�b7=���$���(ԮR�J�(�rP�]�O�%϶#�C�%���z�އܸ7>�����>8e�l�R햠��_䵵�p`��.!(��Q\+O���>���P�)'��q[.s��)g{���C��� ڀjk���r4^��Q�����ed��Cvm�=����6�;X����d��ok}��V���ܙ�.+�=�%�ƭ%\势���qEu�����%�l6�ʁV�ܬg�_��&��"�&Ev��Gn��i�"�I��Co"�Jg͑��2�
N����*J��ԞRxI��W�W��O	8Ωg��`V0*���>��I�a��l�07��BsqH�R'��"qH�R'��"nI��f䙹&nI��f䙹&rH��_�f�rY�,�2'��&rI��&���f��B��-���T�!YVB���g���I[�H[���n����Y��
n�B�b�X�����g�c;�����Z��
�RpD���C8�oE�ܡ�֬����|K%z��-�I���-�Ȼ�\	&���ʥ����K�s��\��,�N�*��R�N�*��R�N�)ԥR�I���4�&��+�eR��U��dw���6G���3��|3�ϋ}�Qo�J-�k�wd��vHwf�ni���E��5�����[#�P�Gܢ�+�1]�K�@\�~�J��+8d
Gv����)��qHW-�!\��t�R�1HoH�!�e�P*����.P|t^���A��z�������Ǐ�?�ӨYmӨYm厖��-c�:Z�C���C���C��ޝt��:�d:�dX�^X�^X�^X�^X�d.X�d.X�d.X�d.X�d.X�d.����Ix�Ix�IB�C��d��],��,��˧P�˧],��P���,��],��Rӟ%�5J�~;%\t���+x1�ӟ%P\u6���n����t��t��t��t��t��t����.���/,x�C��,q�C��C��C��C��C��Aq�Z�㬵��U��U��U��U��]#������M�,�A�,�A�,�A�,�A�,�B�,�B���.☸#�#�8��l�R�J�/8�E�M3����j|o��q�(���|hY����P�l�x~���`ˣ�T/L�y-Z�Z�Pmw��*u��?�=�^It!�g�|i�{�����Ԡ!��M-o !�}�&�}��>�K[�8<i8<i8<n��R�K�sӯT����:��5���[�*��%lw�r�D�q�H+5���г�!gw��vr8�HSS�춟#��|���2_+�|�[�䡙)E�>B�����A��l��Sd������>�t3�C>�l3��>�l3��>�l3����~��/+�!�����G�~4^W�E�~4^I��d��6I��e:]I��d��6I��e:]S��%:]��P��
.B�¨T�U��d��Y ���lF���v�j]��lF���v�j]��lF����|p�>8c�1ώ��s�9��(������sߔn{��~Q���7=�F�-C��v��ߖ����;~Z�o�P��j���rp`�'���rp`�'�-C�%�$�䖡���?�Z��KP��j���rp`���Q�rJ1NF)�(�8e�r��o�!��˞ܵsۖ�{r��nZ���>8c�2�?�Q���7=�]�o���������e��*9s�|p�j]��K����R�P�S��P�|�$���s�R�bď��t*I�)ҏ�B�G��v��q���^/~���헇�u��U%Sa�R����}�^��Q4��EQ���#���5�P�܌qF�#��K��%�'����,����]�[���S�u��4�%��vO�*�݉`�RhX�iI�Y�ړF�����}�}%�FD�>������H�3���c	v���<L������i?�c��K�>o��持Au�ۋ�9�����"qH�R'��"qH�R&䙹&nI��f䙹&nI��g$��I��nK7%����"pț�&���f�~Y�,Ьn�Ϳ���o�8pg�*~`��T�vK�5��5��5��5�k�X׾��};r�;������ŷIN�HZ�Krzm�򺬮�+��d3���j�e��wz�j��vŲ�!$���?�_k*���dC>��"S��� ��KK�RՖ�zT(>}
��$���T��>�ϡA��P|�N��B��Jt�)Ok�)�ue=����ו����V�gž�(�ݥ !�Y���������>��\Qf��E���d~�X�y"�+��I}�K�@\�~�J��+8d
Gv��R�qHWH�"#8�t��!Y�^���gz��#��G����?��?P�<N�e�N�e�N�e�N�e��:Z�,t��X�ksP)�sP)�%�V�K���ǁ[劁 ��@�yb�H:s�Yt��������Jb�Jb����������b��b��b��b��b�祔��2Pg��(3�̔�YJ�,��=,��5�5�5�,��,��],��Rӟ%x1��/-�PcSP~>V��A��+N�d�\�P\u�N�Y�*/�<	N|	N|	N|	N|	Nj.��0�˧0�˧>>/N||^�x��:��zu���������>;P|v.���]A�2�qҔqҔqҗ-�,����yoe����^[�Yyo��.☸�b�,��*))x�ĥx��2^6q��DX�4�c8�x��,q�ȱ�k!o���vҡt����@^�� ^^@��O�q�4tyN���#�J�(6�P~*�A��:sܶrǪ=�>����%ô���3�s�3�K�3�K�3�K�3�K�.�/Nz}9�A�c�Rӟ?N�P:��*�Q�?O��6�[\۹o/O�]2�x27��d��@��ޗ/x��Y㵺��qM�[#��̬��	Y���M�|����W%߮%f����R�Sexb�����M�a��[V�u:�S��u��[a�u��[a�u��[{�������_y��#�/+��/$�a�N�$�a��.�$�a�N�$�a��.�)���.�B��(Px�
�
�R�VH?��d��Dj]��lF���v�j]��lF���v�j]��lF��(������sߔn{��~Q���7=�F�(������sߔn{��~Q���7=�F���rp`�'���rp`�'��m��~��߮)��m��~��߮)���m���|v�z���m���|'z��m��~��߮)��o�������)���v�1NF�(ö�0�>���m�a�~�'������n|2���-A��_'���-|v�>8c�-���Q�v� �����̫8�g��=�;�I�E�i/m��rG7��6=�k��������ؼ���ɜ�K]-G;$Si6�w}�?g�dj�+?f��`d�1}޼Vv�PI?�De��F��ԟ2"�&��ݳ��_V'V��;���7W��K_�������o�zH�Wړ�F�iI�J�mF�� T��jJ��=��D��O�aϯ͑_q��p\ѐ(������*O��@� Q�(�OT��4&�&gۋ�9����)�D�8�N)�D�8�M�3rLܓ7$��3rLܓ7$˔��������f�rY�,ܖn�n�ۀ��v�?%O�S���g>�9��������%W�ȝ�'��,rI����!�8V�̊?�0/ߓ?$J���8�H^�Z��f�dK.J�l�n鴙Jsݰ���/�햩w(��w��݆a����^�j���R�/>�KȡR�%:^�
��)���T�*/^�KסR��T�z/^#Kה���M�e��B�nж��.6�y���k�����1���ϻv-�7"�cr@~���O�ri��N��ߋ2?�⽰�K��\��<5
Vv���帤+�␮��CzF)�,�/Y�^���Agڂ�-��[j��Tm�?�P~=:��zuC���C���C��ޝt��:�i�u��yb�H<�P$X���]9�,�s�Yt����ρ!rǁ!i������ρ(t���JJ]%%.���IA�K��ĕ�PbJ�(1%t���JI]%$�3�X3�X3�T�	*��x1)A�J]%%(3�9.�����-:�2\��ezK��t���@C�� &�e�������T��劁�Ӫ���~�%�bJӨ1(i��4���4���4���4���4���:K��:K���K���K���K���bJ�%:�e:�e
���
���
���U����T���.:J�>K�p2H�d.���]#���G(t�P�.P�.P���.☿8��l�R�I*�X�e|l�+�g���i������:�[��b�ʋ<*���;�4,�T*���Pc/ ^���5�����T)-��Tze���Wj��?��P�ʎ�B���P�K�ӟT��8wI@p�ܱô�� ӯT��qM:�G��l�?N���H�d:�+i���T.���x27��d��@�E�Y��0�ax��ldq��dw*���fVgd��H	Y��d�W���P̏���ġ�^��A��l���0ă��M�������+��ҿ��+��Ҽ1m��l�[exb�$���O�?)�"��/��G�~4^W�E�~4^I��d��6I��e:]I��d��6I��e:]S��%:]��P��
.d��Y ��H?�F���v�j]�ώ��s�9����|p�>8c�1ώ��~#s߈���7=�F�(����ᖡ���;~Z�o�P��j�-C��p��\?���C�;��N�;����C�;��N�;���t�.�R�ӊ\�qK�N)r��.]8�ˡ �t��]wN�Їqt��]˧�t�^�)r��.^����xb�/{���pcЮ�� ���980��;�����6��?�������\oȎ�#��z�7寎��K~�R߈��e�?o��@�T�<��O��Ӱ����:���rE��~�ƠG?R��a�)H�F.7���*~�{n��N��
�;%l-�;8W��C��}(�>�b�F��PXѷ8ʺV8�,3dBN�
U��"�J�%�T�d�Wct;%�5d�i.p�-4�܌xVp��ѿm�w��Y���K����-"t$�R(՝��k"Y����rȚ0Z9�Q�7�sýƁ����q���sAu�ۇ�9��?�@�}��E��O�i�H�R'��"qH�R'��"nI��f䙹&nI��f䙹&\�WܤWܬ�+7%����f�~`���3�����0g�*~J��*�p�9�0/�`_����v��w�X�`_ϗ��a����eTb�a������1�Q�P��4�1��U�,��[V�U�l�셯/(na��Ѳ�NB�i���%��[o�e�Ҷ=��½���1�d�rI;˗y��b�6D3���ix2�/J�KסR��T�x�/^#K׈��"0~�%/v�KݲR�h[]��r#�ܔ��R��W�vw����1���ϻv-�7"�cr-�7$�O�ri��N��ߋ2?�⽰�텸�o��¼iY� R�!edC����b��2�"��8���)�����oH�-��V ˁ�TN�.:�P�P}-n��e6��Zޝt�C�
o,T.�x,T.�x��,A�.����2IA�^���^���^���^���_IA�K��ĥ%%%%+++++++�^W��ĕJ�(1%t���JJ]%%.X�e.�ty^���9�r�u��zK��A�V�d�;���Է�'�^�N���@Ώc g/��?/ʐ2Kk*IU$�X�W,x2�,A�+�<K� ĕ�PbR厖B厖B�.�B厖B�Y(i�K(i�K(i�K(i�,��JU$����UA��*��d�P�J�(Y%t�B���8�p2H�e���������,�P�K��%(�e`.q����W��2�6q����",ph��i��������[�k<hY���.���}���_aP��^@��N@��O��dh���9o/O�ͺ���TA�A�~���������=�=9�G��Ӟ�z���ʃ��u����/Q�?N���-�Ҫ������tt����ǃ��Qz\�Y���z:.g����w�f�����s���M %f����]�VJ�d|�߮%f����R�Sd�un�$f�{��o�M����_�N����_�N��l�[exb�+��'��}��Oy���~��?+��/+��N�$�a�N�)��N�$�a�N�)���.�)��(<B��Y ��H?��d��Dj]��ls�9����|p�>8c�1ώ��s�9�����n{���F�(�������a�2�;~Z�o�P��\?~Z�o�����wo��އrw�ܝ�w'z�އrw�ܝ�w'z�ӊ\�qK�N)r��.]8�˧�t�.�S�������p�.�?�������p�Nr��8�0/TR��\�QK��)r�E.^��'z)
�E!\���rp`�'z��r|��?��R����R���(����ߖ�8c�-��K~#��Կ=_��6�e��d�h{Ij���)K��!RzuIY���T���)H��Hn��Xܟ�%r�����j��k918�����=�e�՜b�%�VEF��g���D�Yϲ��l�n�7�o6~����7�	M�f��>=($��YȤ��̄��	�D�7�'�O	j�7�M~m�y4���q=P��k7�de\
L�m%Q�� g�Nh��c��p�p��G��&���9�9������}�vE��O�i��Q�ȣ�*��*�Ƀ~��Vk��~Uwo|R&䙹&qH�xߕ]����gv�f�7$��2�&\�˔��"rY���U���+��Wm��c�b���hT��,v�9�,�
��*�p�9¬�
��+
�B�T���һmգmգ@�!��z?��ꭺ��귺�멽�/c��\��F���$��~��%y/X�^!+�7(_=�^Ej�~%T*^���܆a����)�{"5-(��E���7<�j*��'E���5-)F������������2_��xdq��.����.Ql1ɧ�=��8��Y�:)��H�څ�E�q�,R/P�H�-�#��G�nq�,�?P�<�P~<��P�˧],��5��=,��P��P���Pu�P~<��<zޝt�,x2�<�"��� g%i�)A���i�)H��]%��Zu%X�e(3��^�Jܴ2[S�i[��?G�ӟ+ r�H��K��i�@��JZv�ܨ	|Z�9��9|�I���@ܖ��C\�t���@C\�`!�t�g�q=:�9��g��ip��Nz<�Gk��ʼV�Wz���`:F��I+����>K�b;_Α��t�����r������t�/��?J�.�P�?���?���2e`���zJIZu�d��JUP%*��rZuP$�9����Z��$���*��*��$���rU%(2�e.�%[�J\����������%T.J�\�x��2�6)%E�RJ����g_8����s�DX�2�7���������гgx�lY㵰����г�P���x�����rގ� \��R���$�?�IjH��ڃ��pe�u������
��]�(6�P^��A��u���]�̷ R��P�m>�����<oF���2p����^?�@q�ط���<�-�6P̎�C2;�ߕ��fVg{�Κ-�qns���~JW��(fG�]��P�d|���
�,��qe�a��$f�{��o�M����_�N����_�N����_�N�w��'��}��Oy���y_����y'k�v��N�@��t	N�@��t	'k�v��N�@��t	N�@�A�(<B��P��
!B��,�(U��
��~D~?"?��ȏ��G��9s�\�c�>�F�(��evܣ��ö�0��� ���980O\;��A��ǹ=p���o�Q��@;e��lܒa�l��C��w>}G_���Et�1K��)r��.P{��q@q�/U�r�n�!�^�����*�P�=V�Sv�n�a۞��g{�o���������}���Q��Ǹ�4>N�WrQ��I0x�N��Ӡ��>8`;f���W1\��S�����]
�%
������~���(��d�b���a�j���9V��6L��]�B�H�$;[&��߾�M��	KS�VA�)q�^s �J�k��$�nF���#�[ն�hωk�۲iy7Մ
Y�����o����)��*�g�O"1*�Y�$�R���_Ȍ��,��&��9U}�6��������v��γ��8-�h�e��'���%�U�JHDg�d
2p��X\,y�nnnnnnnn�ѿ��s@�Au���(Nk�O:/����{�򫼘7�`߷�;���f�90o�����&nI�R&��0o����*��j�kڈk��ϫ��;���f�rY���3�J��d!Y�E�E�}�}�}�}�}�}Vg8U��l�
��m��Vs�`!Xn
/���"�������o�d(n�/������bۺ��ڳ�k�}�.�R�4ܓ�p��{�	��w#��~@g6�?�i�?~,��>G��;˕
�d���;]ȷ������>G��>3�6쯼܈Դ��6�X����#�|�۔���N6���ղm{$�6짼�����xb��J�-��VP"Ď��,R/P�lq�����8��\�?�xmB�-�#��r�:�P\u7�x��X����l�e��58�����x��y
��YB���:9+N|�C�2�,A�+N���Iq��X��X�UC�2�,A�+N���Iq������d���߼��͟,�͜�͜���@���5s��4��t�/��a����+/�� s��Ӟ?S��t���r�����Ӭ�<��i���R�>?%���2[M�\�V,p4�fK�e?�C���r��eXcY���I�g��Voc8m�@���)'�=������[���;";�WE�H2��U��`�����ӽ�5sʐ3�����i�@��������t�/��5sʀ����._- \t�P�-A�WIr�m:�q����?K��~�%PU%],��<|�-�.[�����%T.J�\�P�*�X�eb�)%E�RJ��#��2��8�B��3����j|n;e�q�(���bǏ��v���ر��<hY��f���~[��j�#H��.?)�z:gH��2���[+kPe%��e%��e%��e%��#�J�̷_�|~��e���ݿ�W2܁J�UB�����"�L�~R,A��X�rqb�j!oK��g�@q��g���<��ܨfGr��Yߕ��fVg{�Κ��XfK�ey���~J��~��"�!C5Ŗ�,��qe�a��$�����S{��l������t��J��t��J��t���I>������{ȼ�����h�����;Xl����t��K�Jt�
�v��N�@��t	N�@�A�(<B��Y*P�!B��,�(U��
��~D~?"?��ȏ��G��9s�\�c�>�F�(��e�۔a�|v����rp`�'z����xcܝ8��z�Ѐv�qN��� ���x�<+�A���.]w'������(=����q@q�(=��nz����f�·����v���{�� ��C���(=���t!�}��o���z�������-��\_�SݡAΆgz��)��zv��k����\�!xΥ
����{k���ߒd}c׵�J>迪)r�{��)%Dd|����D��%�G-���u��]���4��oġ�����y+���cS���Y9�dЍ�c?�*�N҂ܤ�&��X�"��2폔�"�9%��)<
E�g�r(��Ԫ%��A%��?��,�I��Q7�K0�K0��]�@�y�y��_������u��q�g	�����\,`U�R�g��l"�
��F\,.��7���������n�s@�}�y��.����.(��W΋��'Ł=�6�vDݑ7dM���,۲&쉹f�����,�:V��+�o�o����<R'l���U�83������.�+!
�D3�@Ҿ��|7V�_^�_^�+!
�_
�_�*�*��U|*U}T�Y���ۂ�J�܅�"q����z����辺���)��ƒ���jη�|��FP�Q��яȜ��vP���lx
e�sS��R�QnsN��^W�p�){��Ƭ���k�*Z��Y_k�q^س��Jt�*?���p�G��t�)%�;�?~�9%z�~-�8b�/�s��Y�!�6)���~,H�E+!��VCb̎��ؤ~,gފK�4��$t_��+#Ǧ��K(r���������!A�K(rǁ��<����vR<[83>���������gIr�nX���{(|[M;A�N��u5����t��||_-��C����r�n�W<� �UAT��.�9��x�=��+g��W�t�O֦����E7`ʠb9o)C5�c�q�V��;ޒ���[P%	&��z���ZC����H����--���?�;�V{z��{\�]�+����.x��J�P� ���%	�dv���P�I��a�{�<v&2Iz�[��T�ez��qK-Axi+��I�{=9��]#����.��\�����{({-9��P2]"J"J�i��b*�b*����,��G���.:J�\J@�쬁q�Y�t���@^�g_8�x��"���b<l�+�gX��i�n;8�g��l��)��<�������xг��BϔX������_aj��x��9�:���d������oGL�2@�y"@�y#����-��������^��%m*�r����U�� /�L��R,A��-�2~7���Qz\�E=��ż��v=�i��W~Vk;�Y+�:��s���:hfK�a�/���~JW��.�q(w�B-��3\Ya����Xf����/�M������+�+r��+�+r���+���N�$�+N�)񭲞�/)�"�-�~���ж��%./d��씸�F���J\^�K��)qx���c�*r�@�T��<*9�G �F��(Կ%���k�Z�햾;e���k㷃s����x7>\?���ö�0��� ��C�;��N��� ����^l���"�J���|1HWr��ܶ\�0�O����[.^ʎ�B���m���}�e˹l�w-�/}��C�������^�*���}q����C��G�<4>��U����ܫ�]���6�0�}v��z����/�ܣ�*r[���{;�j�+�)�����)����t�o�ٷ����8ls�[�g2��kX�q5�C�H�gύ���5�\9�[}r�
H�}�(�*�I#�8�=2!)n12��cK���^үJ��)5�"zPWl��ЉdJMFOv6_�,�|����)g������"�Y�$PI7�|"���ʿ��'����^�����0(�o���w�;�]n�u��q�h��w�;�n�(�'�'�o�O�$
p�3�q|M�2��p�p�p�p�p�p�p�p���v����s�Ђ�V'��O�xN�wdM�vD�;$��3�L�8�'�fܳnY�,ۖm�7��.����h����r@��4p�Q�Y���Yx��XV}�U�83��o��[x-���*pʜ2�nC�>���ϟ�|�2.�g��"�7"t4^�X�G���_��?�|_"q|��s���7I�E��}ucI[�V4��%�V�ƽ���/r���w%���2�M��� Ճ�lx�~�k��|��$��Yd��C8�^@b�ދ9�ж�R�ƭk�q_ȳ%�{�m��r,�}���Ų_�-���9�i�!��ȇE#���E��+O�hfGE�n�xt�i������oNy|��r�^X�䪃��$���d���2Pe2U��􊁒�<������i�G��,����\�<1M�O��I�v�7r���j�(:PmvE��)y�;=�u��_����x���s�Ǌ�p�+�mJ��R�Y�Լ
do���\�r/eG#8������4�~�@�Ag�W[���|gP}Ky��op��i/�"�RًT쨤�:�[D+�%s�d�[%,4B�R����p�$���v"�+F=��=�������n�}�Z�[ϲ{����zJ������ӷ���||�C�9hk��?����yڇ�]:�qs��t�gt�gj��T@�T@�TK��>W���^[��9o���.M \��p:h�b /�����p:j���/�񳌬-�1c��B�S8�f�#��g�E�;[P�_D�}�c��E�{��8[=�z"�,�x�.^�D������&������+1bV|oF��4��� /�Z�đ�A��X�$h[P+1f�bz.�Q�T�Y���6,�i�?v-�u�����I_8�w�f��+5��s��d�ZW���^K�;�����d�&�����R���~��!����^��A��������Y{��l������ܯ���<jt�ƧI;�ē��I;�ē��J|kl�ƶи��B���[X����R��J\^#��`�،��b0xlF�T�ʕ9R�J?	G�!(Կ%��R���;e���k㷃s����x7>χ�s����}p��\?���C�=p��r��6���o� ���7�8���ÿ 8��@�o)�5o��{�=8w�r�r����8�������a�>��'r�r�[.^������B��^��ܨ�w*:�:熃������ʎ����ܨ�A��ߥӇ~xa��߯��xa�d{�V�]�}�C��P��M�^��ӊp�>����bdܼR%��t�V����E(|Wn#�r��k_'m�� ��5a��̽n2Aң
�]ۖ]ȍgء����x�K��D��a�]τI��&���'`D��e�_o��9TM��<������7���,��'�vY�,����"&���ɿ�M������RuRyXyW�Y��>6��6����_n/�q���:݂�v��`o�����N�`�݂�8�d
2�q07�@���N�~�_��p�扸}�}�}�}�}�}�}�D��c�^&�Nh��`���� ��Ac��������,k���d��&vI��f���w�Y�Łw�����w�Y�Łv�G�"���政n}]�Uݼ	�w1�7mCu��5e�Y�2.��8eN�*<��w�/�Oor�qY��ߙ��ϟ�|�4�����D3�Ȝ7�G���4^�����{;���Tb�1yUؼ��_"q|��eHnB���筹nBې�i_[ջMף(qK�W*�U�����-&#u��[�X��(�1-��jܭ���4=Ά�!��
�E쟨l3%��8��Y�~��ێR�%8cnZ���xےL1�Ⱝ?9�i��@Ix�[�¡l��T.A�*�)r���?P~J@��/��V��qN�ed~I�!^����l�����>���D�u�	-!ɡz�D/A���r.;	��U��N6Z�:JG��f-Rʠ�iԲ�����d��)zi����jh�Ta��;*�d���T��7*��i/ţط�!R�N)(.yV�Y����;$�IH~U�)|�0Ʒs����8O��EKY/ �ݡ�
����h�mS�ݨ����,t9KGV�!Q��Ua�����-�����b1ǲV��+W<���[�NB����))K�y]z\���
�#Nd�v^�&�[[�||�H��Zs��d~�|����u��Nx�O,x9nX�r�u3�P3�P3�e��˥�t�Y��>"@���q�څ��j��\v�i㳵��@^�gX[�b"���O��jb���H�L-�vpw|n��|}�E�kd)����E�oz.;{|~�-��������K��af�,�̈́-�r��şQ|DY���P11c��Ŏ�'af&��LY��~���t^>â����v�@q�ط���<ǿ�m%|�e+�)_9���ΦI��i&K�y/��q\��#�R���I5ĥ$��������\3\Y{�����{��W�Yeu�I�H2N�A�}չOyN����OyN����OyN�q��.5��ƶ�6��&�?d��씸����R��J\^#��`�،�P#�*r�@�T�ʕQ��J?	j�
��p�G�!-\�R��-\�\�����z�ݼ���v��ݽ�z�ހp��ܝˡ �t }�B�Ӏm����l��@!]�g���\i�D9{}˹�piq�eGv�o��!^�����r|��}�e˹l�{�|^�����w!z�/A܀휞'�=��9!z�ߦ߹�ܻ���e��S�z���M���Gt��1!p5��nR���pb[���$.�R����@u*o�M���JV"&��ȷ쥖�;M��l5w��Ύ�%l)��r�o!N�d��JW+����JU��c}���d�ÑG"��ȉ�����}�=���%��|m[8��XݕI��"VR4i:ѱ��'�FY��4
E�*���I/"�9g���'I���F��:�|�7ʿ�Y����
��b`o�q���:݄��O����$�|�&�.���8.���8.���8.������Y�u�ۇޯ�PW�����������������*�v9����Y�����[�t�8ba(��~���'k���d��&vI��)�ȧ�gۖ�,��w�ȧŁwr����L�.VnL��Wh���h��*���?�{r2�v�+v�潮Z�9�y%S��o�3�ϜC=�D3��7=�P0Tt	�0/�`_@����|"�^UF/*��]�ʐ�R���`����N*CeH��m�V���Y�{.�[�r\Te�캪�B�*H9m{-���xk�����<��+Y�x�������d{n�nJuŶ-��s����aZ|��E���P���H�l�eP$.���zGKe���!f/�����V��!��B�Y/n��5�a�9���lh�r�~! �<Z�%!�UK��}2�T��|���h�b�I��,E����>���*����C�HvI �	I��I)����l��vUjZ��2ӹ�W<��\�b-Mߌ���3y����a���ͦ:^��ej�����nǤ�PT�%����vʩ�S��Uc�+P	+�qA��T�Z*2�8�/�B�]�Ѡ�V��l�9
�P���Xh2���/P� �@���a�m�Ke �\P�v��+T�OY/��rȏ��||�p�^oVO�_�������L���c�]���=f����9��555�e�
�gj
�gzD,�t�Y��>[���i���e���\w���i㳵��@^s�D-�1c8�E��- %f���2�ʅ��,��ދ������@b��l����oE�oz.;{|~�E=,�i�w�O�Z��l����?��i�/��̿E�e�.;/�q�}?��i�w�O㽺��-�u����x�8�����W�6RN)ʒqNT�%��L��Jx�vS�s�N+���|�+����\JRMq)J�BW�b��/���{�����exb�$�$'y �;�I�H2��)�)Ҟ�B�V%=�:�ƬP����d���X��k����J\^�K��)qx���c�*r�@�T�ʕQ��J?	G�!-\�R��-\�R��-\�R�����pa���wo���v��ݾ�wo��ހp��=�B)�Њo� }�Br�@6�p��n�m�p��S��A��@!P����s�����Q'�wi=�HW����>w�K��-�/�{o�l�|��8��r�r�[.]�e��C������>(^���p���^ʎ�O���D*?W����������u|zgO앒6G��[��l�d&[���m�6���;#��REc,���YN��vA���c�.T��F[og�-�{!Vn3~X�sqX;p0�D�P-*I����X�cZ�v���Uz��,�Y�5�0�XUҍjض���RU�}�|"E���j�
��k�j��Փy�"��E��g��^��m�M��O(�d
7�7�7��?��Ro�7�|"���07�u�	��$�|�7ʓ��c�����8.���w���n/��|oZ1�g�q�(�����(N�����������������4m�T��MjO/gc�Y���6Մn8�)�o����{V��'k�ݒ��ɯݓ_�"��,���+:7,
�,
�Vtwd��K'Łwr���vD�6�'�*�ÑG�>�}��U����pg����rY�Z�4��3�v�Յg��Ȼ��v*���J��!�Cr܅=�~j�HVz��d!Y�
?�|>�nB?*G�yR/*D0Q�������0U��7= �2\Te�캪nz����_!na��1�:��M�<����j�[�~����,�NT$W%�����?%|�M�.[P2PǦ��:/+���'��9ƹG8ܑ��B���4�U9G��r�d~Ʈ�:���}K�R��-ck��K�Q�l��vU[;[]�X>v�U���@2�~"p���J@2S�eP�*�~"u,��v�?+v�C����T:J���FBTe%JE4�~�w=e��?�;]���!����1��XjZ�{�Z�NBPqj����
����
섐�Um��J�R�S����)z�j�!Z��2�<GZ�V⧒�S�f��Td�+EG+������r���?a�o��7ߍ4OƦ6�)@����7۞Z&�����s��\�\l�ew���]d��&ϧ�Y g��Ӵ������A���A���t�G�ӯYP�cSP�cYP~��\�t��[��o���>�@�촁q�i�ܷ��r�Y��\���8�x��"�ر�e����L���5:~q�賍�Y�6:~q���[�m"�i 8���l�.;{�q��?����?v-�u����� 8D[�������)��$��oE�|�.��p.���H� 8G8��󍌯�l�|�e$✩'�Jx�ZS�2�L��I2_-)����Jr>J��|�$���\JR��P��R�����0ą��H=�ԃ+��^��;�I�H2N�A����OyN�����B�V(\j��X�q��M�~ɵ��6���./��씸������<6#��*T�J��P%�����~"��-\�\�����pa�����v��ݾ�woz�ހp��=�z�Њo�"����N=�ӊ\�1K����\�1K��=��rz���������܀B�Q��|>�[�)U�����~+f܎�D��˗k��/��C��E9;�NO|{o���Ƕ�{e��\�{e��C�B�J)#dg8�C�p2F��e��ɫ�uc��M�l����>^Eo���$�č�����$��}�j\R�ؽ�+n�^���o����Y:��_<���F�_[�ё�O>�'�հ��9TbYװ��c|�,�jɮ�K/��I�'a�,�ω��~�c���gFE�&�K ��Ĳ1�ω���^E֭����(���^Ź&��a~l�gc���a��H����"M�"��W�RyF�p�3��RXK!�E���'�d
3��y������}�UU�
��2����������FڕI�$T���2�$Ѷ�a.��mRD��v���V��^ד�%��OvM~����d�{�k����������Y�ݓ_�&q`]���r��nUw�"�E�����nX�nDۑ6�M��&\�˕��"�n��ݝ��eWaR��h���T�ʐ�R*Cr�]
�B�ߚ�����d(����S����B/���(���n_��3�`��c=M�Ss�]V/�x�ʸ�ʶ]�zn�Zޭn�oe�r�B�FR�P�Yt��KU��i�mV�mO���5�1QߡJ�_y
�jr�������Զ�gR�jT���% �)*X�/S~�eV�@4Ȧ!ʭ�R=�[%%�RP��RG�H���eP�C����*�~V�?+v%_��II����U��nò�Jp	) ����+8~"p2�\���r���7a���2�fIK�Z��k}m�K�$���U�RC���<Z�(_Q���rThrUX�#SMj)��S�ݨ��r��/S����8�v�5vP�J��ұr���:W��M�٦���y�e,���;;��� �}�ea X(�2穱�ji!�h�v&�����i���w�(J�#41����iσ��;�-���t{���=%��4��r���?��^*��Ʋ��Ʋ�\�t��2�s�#��t�-�<|�-㳼�����,���-P�4�4�6q��D-�3����X�Z@b�h�Ge����;��-?8�Ş{ 3����6�����E�kz.;{|~���b�[�:ط���;{ 8D[;�����~R��t\ˢ�>]��D��}��J���W�6�N)ʒqNT��r�9���L��#�Ҟ+���\쯊�d����|�$��RMq)J�BS�J��P��X�&���ą��H2�1M��l���d��$�$O�M�����B�V(\j��X�q�.5�ɵ��6��&�?���4��F��A��<^9��5(l�R�J5(l�R�K_	k�!-\�R�����pa������B�0�W���~z���z�ހp��=�B)�Њo�"��8�'N=��rxb�/T���z��/TS����G�����|S��D=1��L���p5��N�������ύgY[�t ���o���/����G��x�o����p���OݳnKP�|_�_vE]�@ǹT�ܯ��6����KA�w���#J_�{�G"A�z$�L_%�7=��e3�[q*n�^�%"�}�Uc9U}��81�e�)V|JU��j�ݰ�J�(�ɹ��;+�dF]װ��avU��`F�,o�RNOH�F_�G>2_������[�����dщg�c"
��2(�~hȠo�@�^XZ�7�H���ՕRQ�A_c��각���� ga�&��B+�� Q�*O��@��Q�VR�d"Y��W�W�RRyFu�O;�tN'�í�=U�U�T�Q�(��'�'�'�'�'�'�'�'�Mk���6�|[;���4�﯉�/���n�*��{J��'���z�v���,�d���5��+��x�h�`�ەUݑN�f���&��7��N�f�7�Wy0o������n}^����7ܬےf䙷"mțr'%����f�n���Cq�%W�%Hn���y�5T)�s���!@�P%HnB/��硹
�
�~Y�����ʑ|�_=m�G���;=[�V���Y�:��u��u��:��:��=�.��}���-��[���W+ri��n&wm��r����U��V��Y�y����K��M�Y��n���J�Y�-�R��T�%R�R�R�R�R��R��R[%$J@$�?$���)��R% )ǲS�IH���IH��IH�����������>1>!�\�vY�_�_s�Q��ò��촼SV=��l���rW�e)��O��J�.�VP��(�e
59J�NR�S����*�9J^�)K��QYKFP���T�Z*y-+�FJ�Q���d�t��+qA��hx���G�f#�{M	�}�i���h(��
)���e�!�h�vZ2���e�.yh��Z&����y�d� W?v�&V�,��J����N�,L��N_���ˤ�}��z�9���&�ލ;~��P2�5�������r�M9�u���G���;%P��7H�59]"k*���3#�.��i�ƧO�5�nq����-�628������O�B��is��E�m$q����-�6�o��x�[�m"�i����s��8���Ml��ob�� 8D��}o݆s��8��r��)��T�+9RNs��ef�I���O9�I2_-)��*W�$�^���z�J�Y.��%+���JR��P��R��b�bB�a�
S�Ye?u�S�Ye?u�S�Yh^���[�{�vM�:ɼ�Y7��&�?d���X�F��R��<6#K�G ��j��P8?���!ӀD%�<^Z�[}Q����!޹�878��
���;����;����G����t#��RЀv� �o�
�P��1��k�Ѐv��{~'�=����8?���vz�_���$��g���*�r��(�=�������D)�_;�D�� ��7��I9̡�ҳ�^�߲+r�r�i_9��t�/�'�d��j̋��Ӹ�u�VR�.��J3-Ħ�61~��n��vu�$C�"mɛx�S!�&k��v읹`�vW�lU�����1*�J��ύ�c1*�J����`���g�D߃<�8D��E�&��}H�/�A_"�<���s�h��N�&�Y�_�v�&r�D��E�"���v3����NM~mYU���r(��(��x+������F�F\#:�:�:�:�:�.����oTl
��������6��F@�:�3��:�3��.<�<�Z<�=Q�(�3��F&�No��>�#ѱ�/a���,6?e�~����������?zՄ�w>��`ϰiW���U�Y;VNזO^Y>�5��+��w0.�`������=�	��Oo{x������'�*�Ƀ~���W{s����ߕ]�����"mțr'%����f�v�϶�}�s�������7h��W�4�Ҝ_Jq})���Ҝ_J�o�4+�Cr|�Jq�)�0P�R*CeHnB���!�
�|��i)ڳ�u�u��]��]�u�u�{bB�b�'��/�x�ԡ�9Krr���\W丯�q1mg#g��Cg$V���*���6���ڃ�-2��\�Ȧ���)�� �K��W��W��W��W�$��I*�V�?+v��JC�H~I���)����%#�)Ǥ�zJ@$�J@$�J|b��!�|bd�� �;,�gg�_�U���4�����WzJ���Uh9*5J�NP�+���;|�F�(U��k���vR���R�\��KvP�]�-Ee,qYKO%����S�h��Td�u+�+qA��Pd�W�+懕��BG�Б�Gئ�
)���gb`ؘv&���e�!�h�vZ2���e�.yh��Z'y����T�=7�vW�KS�G�%�vSW��\�{g�[+2]&�V`%��P�u��*
�l�m:D,�����<����G��>�M�8�*��]6���W-�4���\S;�b��8�x�v�qܨ6R�HS-�ȷ8�C9��-�6=��c 1M�-�6>6)��M�-�6�q����@gH���E��-�6�o��x�[�m"�i�H�8���;g$��_�����[�wa��{��62�)���g*S���^Vr���Y$��L���<�-$�|��\IR�q%C5ĕ+�W���Y)^��8bR��R����$�cB�1rL1!Y!�,���!�-���!�-y нջ&�d�S���u�yN�mm�M�~#K��iqx�./��b0xlr�ԡ���C�/ӹ�|0��m���:!޹�;�8�B
�C�^��z�އv��ߝ�C��t#�R!ЊB�0ބ�� ��G��v�O��s�t!�;��@qN^�r��/M�v����*;��r�������-��)[�n���ؾ���H���c�b�[��؈^���;||����q85�u:���ҿ+�o��-��~uE�/�n�H����Vjn{�N�g�Y���rK��#��'iI��y���^үg��>�y�3ϱ�}��)��K%��F%Q��JU�F%Q7��N�g���՜"E�"���`}��pWȾ�E�vpW��Q���g|��M���&����?���Y�t�T�V?����|�2��&rx+�x+��o�����'�l
6p��F\#.�˄e�2�p��F�F�R@Βt�3���gY�u�gY�u�gY�u�gY�u�M����.h��gY�����Y�s�������$%[��?e�~��BU���I	V7���a.(�\Q�����܋E�"ş`ϰg�4��U�Y;^Y=yd�$���߹�ws��;�x�Y�Vm�	�ʮ��Qߕ]������U��)�)~�<�7�H�+5��r�rY�,ܖnK7��g>�9�������0/�J��d!Y�z��8������u��u��s��C�D0P܅�V�we��ƽ[n�ؾD�
��Cr�%cIN՝;Vu�{�z��:��{.�:��:��=�� �$ą����c��7R��Rܜ��9Kq��J]�+���k6ވRH�ݨ�qõ���kW<�~Z�~��!��?L�gP�)���)��<��\�v!�!�T;*�eP��C��vUʢ�TS*�eQL�)�E2��U�N��?8~"p�D��g�Vp�2)�[1�"q�D�؋�LEX�WS+�=��l���$�4<��NR����e벅��J��P�]��범�W%�+�����e,qYKVR�S�h��T�Z*2W:��Σ%s��n(x��<��Wͳ�و�l��b?�4�QM4; ���3�0�d;;����67=M��YIs�R\���=e%KYIR�Rq�5�]���Is�D���a�_��X�W�c	�j+�ڟ'~Ved���#�I�R7,r��;x�=&��:M\��c��T�A�@�T<�T<�i���1�:��尳iP��TX㵑c��B�Y���v�3��q��qMO��9���6Ql��tR�e�J͗E+6RVl���C2�eߑ�)&Gl�|Si+�I_�J���W�6��)��qM�3�m$�Y��ef�W��>�)���_�I2;e$�픯+9R���I2�S$��L���d�/��d�ZI��iNG�R����z�J��|�$��T*�%)��'�P��R���(P�RG�!P�Rr��!�-���w�X��A�����A�o)���6#���v���.�(���.?(����/-A���<^Z���w8oC�/�����p�]�/���_��s�t!�\>�»����;���C�<1HW�)��"�+��z��o���.P?���|�>�*�D=�O�M��l��C�~p�������	O�M��(��l/A����ߊ)e����%G;'��.^��^��;̾�C�tt:{-q%�q���kd�-T�(}��uk2/u�'jm�5���+���
�*Cp+�k���`ձJ�X���"Nϓ�>��c<��R2)�TjUȍ��1���Y�0>�>�`����J�o�D߃<�8D��E�"��H��_�g���
���ϳ��$�W��Q���,�:��<"Y�r(��ϳ������}�'�'�'����$��WdѕdQ���o��}�$��<�<�`Q�(˄e�2�p��F\#.�˄e�7��z�7�� o�������M�&�p��D�"n7.h.o�t>�AsFu�gY����p���?�}�D����o�1�������g��07����w��E�t_*�J�,�E�>��`ϰj�ڲv��z���H��g~��,�:R�9v�'�&nI�x�ȣ��/�*�Ƀ&�9aZ�aZ�{s��ʮ��Oow+5���f�rY��N�D�m��l������3��~J���C=վۯv��F��G��A�Z�vQ���T���S��s�ܳSwp�5h���|�_=�V4��%cIX�S�gN՝7Vt�Y�:��:��=��M�Su�]U�U!v$.�/�(n�ԡ�����J�]��'(k�z�+���z"u��\��W+�����b.ó���N��o5���}2��T����%!�R�C��~��!�d?L�i��D���1�i�D���1�b' �N��?8~"p�D�����b'�N��JP䥳*�eo�IWc�T�zJ��IXc�[V�+�J�C�K�rR�9J�NR�S���e)z�/�a���rXjrU��K5O%����S�f��\�2W:V⃕���n(9[�f�٦��b?ǴБ�4$S;�)�����e�!�h�vZ2����ca��۞��穱��X|k,>9V?��U��*�ʱ��a��/�Le/ec����Z�d1���64�]�d?;qC���2V��ǹ����@�SN���>�f�W9~�6<���A����/g P�Ydv���EAx>���}e��d
�lb���s��~Gd��-�h���C9�[��e������ja�ʋef�-�yQns���<��sʕ�g*S���NVr�|Si+�I_�J���W�6��)��qM�3�m(R_e)�;I&Vley���M��#�R���P��d���$�Y��ef�I���&K夙/���\짊�e9%Jr>J��|�)��*�\d�U�J���,��B���,��B#���?�
#����Ŗ9Yc�Ŗ#���w�X��A�o)���6Q�V�;Z�Gk[�`��FX�`��j��V�j��G�?�>�ީG�w8oN���Vބ:��v�4��B
�C�^�|+���C�;��΄�� ���!^�+� �z���o���p�!�0�S��K���p�-S�A�=�dR�v��;��g�|⟞}�B�w8�Bm����;r�w���-��m��ƌF��W7=O���e���7c���m��om��5=5��&k.Tu�e�T҂E���5��6�ݶhV�^Չd}vX4�Y�D��y��s��ul��R2)�Ԫ5���`�0c1,��Ԋ"��Y�,�L��`��<�8D��Y�@��)7�����PTpbj�>�O���}��&�&���<����g&��Y�u��U��xE��'�'�'����$��We�4l!'c�c�I�I���F�D�D�D�D�D�D�D�D�F\#.�޳��8޳�������M�&�p��D�"n7.o�t!3>�AsD�#:��������n]g|L�07�u�Y�u�ۇۇۋ�sN4�sO�6Dc"1�ύg�4�ZV-+�{V��'vK'�,������;�t���Ww,ݒgd��fە]�җە]�`�r��>�潨Wf>�\;��y0o���o{x�rY��M����f�8dN�9��������p_��+!@Ҿ�v۫F��W%����M��XգϾۥv��V���P����e��[ܗ�vQ�kݬkݬkݶ��۫:v��ڳ�k��ƪ����]��]���A�H=�n�˪�t�bB�H]�^�P�J�Kq)n$��ܗ���������'(n�-Ƨ~{?Ƕ�SQYJ�;-/��ڑ���ͥ�6���*t�b��|gP�B�T�ʖuRΪY�K:��U,��\�us��睝�;;�vp������1�b' �N=��8�"p���"�J�J�J�J�C���䪶�+�%j=%c��V�2U��j�%Z��V��,1\��KVR�����Y�y,�<�j����%h��n(9[�V⃕���:��m����G��w�S;�)�����e��h(v&����ca��۞��穱��X|k,>5��>�O�I��)<e'���}������+�Z�H?*�ʤ��i{+?*������a�����g[I���ey�����t^��ޑ��*�����t��Z�</L�Mg�����24�u�4,��гg<}�-��Z��vv@q���gd��x4[�e���;�n�)���ضVk"�Y��ef��+5��Y���v�S���NGk(X�*��r�X�*��r��S�$✩'�I8�*���(YβS���&Gl��;e+��T�+52L����ΦW�u2L��I9ΚI�tҜ��Jr_)�|E�G�VI%Y1\���Dd|���r��#�ġ�1q��(��)G�!J?�
Z�,��1e�CX����H1�4��H2�֛(�i��֛-R�|=;��z�U�\��V;�(�{��ީG�p��R��!��:�-T���gl/S۔`���:�ЇP:p�N��"�+��xb���� ���;|0�T;����C�{��|�����"����r�@"��?�P<0zܖ�ܻ�Js]ۀ����JA�P��O#c������r�:n��H���kT���M�S~��;/s�������gM�*{)7S��!Z"��@��!gG�Mw"1�^ۑ.R%�L�mɧ�^ױk�]Ҥ�>��+�7s�(�I��I��I�ʣR��c1���`A0 �L$��M�&�yH��_�($�	g;8����E�I���U�*��<
Y�"��
�MY<$������A]�A]��N�_�,�|�
���V0+)<$�|�c��H��F�R@������@Βt�3���������������扸D�"n�g�q�g�pZ'�pZ'�pZ'�pZ'�s!1�1�1��N'�������C��'9����߷�������	�p���C��\n��q��gƳ�Y�*I�X��Z�[��J��^ד�%��OvM~���U[���n�3�Lܳ\�oە]ە]�`߷*���Vَ!���^���������&�x�rY��M�nDۑ8dN�D�m��p��n�T�d"��N/�}c^�c^�cV�cV�o�^�ŎP����e��e��!rf�����f����nV�,4�ʴ�ʲ�v���}7vt���wg�ܫ�ܫ!n_eݜ�ؐ{]U�U!v1{�^����')nNR�d����R�d�.�\Xe.+R���Zn�n���\�^.���\\�rT�z�{��^笗�����Q��Q�jnԵ7Ե7��7���^��Ը��X�k,��T���usήy���gg �N��8�"q�D�؉Ǳc؋�*t*t��9*�J�l���2V��+T<�:���%h��Z(rV�WG+����S�f��T�Y�y,�+EFJ�A���y��hx��<G[f�٦��i�c�hH�����e��ژ�v�&����#!���~�7�c�ʱ��XT�U�.U}K�_�I��)=/i,��%�������R���^�YK���{?�[&�l�]�|�IR�FԵ��^U%/ecs�F����Υ���ez�$��6�����2��{y���X��&Vjc��WO�zu�:K�Zӯ�f�|�B����Ŋ�����v=,��P�S���i�gb�-��g8���M4[#��l��w�f��+5����J�;Y)��d�#��I��H�e�Gk,�;Y)��d�#�����Jr;Yd���s���g*I��.���J�$��L���|�S$�|���餜�M)�|D�%����P�\��G�VI%Y1\���Dd|���r��#�ġ�1q��(��)G�!J?�
Z�,��1e�CX�A�q��A�v��GkM�v��j�[��u�]J��V=u*Ǯ�X�|[{���ŷ�s��!��.�ЇP:p��R����R�;���zp��t���"�+��@q��R�v�`�o��܇v�!ݰ�;����Ԣ�����t7����N��:�y)x���ă��x���Q�u���A�}��?X��;A�H���o!�hz��f��_�#v~=�%��Gl�7���W�B��v��?$�K|>%�&��_k>��*�쉷gwvE=+}#^����Q7�F_�w6�m�۸1�eQ�Tk1���`A0 �L&E�&�yI��_�/�7Ԋ	"�Y��E�}K?��R)?�UT�&�9%�n��XyXyW�K>�,�}�'U��rϷ��'a�c�����v����3��F\#.�ި˄e�2�����������������p��D�#:�3���}����3�g�Ϲ�s>�}̄ƄƄ����q<���3���Ns��8Ns��8Ns��8Ns���C����9�q��u�덥I=*I�ROV��[�loׯ��|��ZV-+�{^N�O�Y=�5��w�Y߹g~���w�Y߹g~��r��,;r��:V�]�(�����r(��Qߕ]���ow+6܉r�6�M�nD�pȝ�s�n�ۂ��v�p]�.�n
��`����ѧvK�<X�{z%Nv�{���|^��*��y��P9.�r��iK�D�âR��(pڔ�����$���/��a�ܰ�W*6^+���bA�Suؽԡ�9Crr���.+�.+�+�J�d��WbJ�I\Te+�-��7r�ow�r͋ⵒ⣈�jv�M�w���S+s�)���+�9B�O+�٦��Z��-\��jZ���M�mKy�o5�c��k]J�mr�>�Ծ2���O�-8~� � dL�b'�N=��{v����%]��Um�Yz���%Z��q���jK�FJ�Q���d�t�:W�+Χ��S�f��Z*2V���΃����n(9[�f#���و�l��i�#�hH�w�S;����e�!���~�6����).z���ƥʯ�r��\��>�O�I�{I/i"��$T��/g�K��R�xm�����q�r.6�E����m��Y���7�9g�g#�X2_a���ɪ[K~�6����{p?^���%J����6T�;�%�9�]��KY#�X-?o�#�Z���H���%�="V�*����-�����!l,�ş-�q��?��H 3���52��8���5=�SS��52Nq��s�L��e�<S-)�iO�J�;-+�촯#�Ҽ��I9βI�u����w�v˿�r�y��ef�I���&K夙/��s�4�%����Jr_$�Y'��$|�d��U�G�VI%Dd|���r��#�ġ�1q��(��)G�!J?�
Z�,��1e�CX��d�Sb;Z�Gk[��kq�]:Z�ӥ��;�R�z�U�]J������-��oB��\��t6Q��|0�l �w�-���^Vl�8|^�P>p
��"�Tz�܊D>vȇ�=
��"�+��xb��T܀B��H�/ �{"�Ŷ��Cax=�����Ԯ��M�V�=�}(6�(o6�u�/�5��nv�j�,S2��?n�#���;/��)7[�B�_*�LW{����[r	R��~�{�X��K�Ȫ��O>2�e~=�?={Y-y3vM~��y����_�w�
�+�`����E�vp���1*�J�1,�K��
xVp����E�"���I�hD���_g"�94"Y�'�I��Y�'�I�Rx��g,�|�����+����Ϸ�yRuXyI�',�|�vT�VU����y��q7.o�\�\�\�\�7��M�&��q�g�3�g�Ϲ�s>�}����pZ'�pZ'���w�\]����4�������O�i��?���4��yƁ���4�4_��޸P6�q��&�������p�/��|&��������4i��\n��T�ձ�V��[��.��]ׯ��|��V-+�{^Nד�%��O^X�7dSܳ�r����$�ycnUV�GnUW�J�Cw�r�!���_7E�;򫼘7��O�Dۑ.Rf܉�"mȜ�n�D�n�}�.���f߳o١X�
�8���n�n�ƭ���B��G��@����gb�q�o=5Κ��@��P.4�x�V���l��iCnԡ�k�VB�Q��/���A�H=�Crr���.+�.+�.+�W+�-��[l�#;��ܙ.+�-��ʵ��zƽ[/;-��.�J�U�r]�p߱��{�;��ܛ�����e1\�:w4;-�������.�5��r��S��mu-����6�dR��_i�e��!�d?L�i�D�؉�1�b'C���䫶̬��J�A��P��rV����)h���d�u+�+qA��P�<E�FJ�Q��Td�+E+qA��Pr�<G[f#���=���i�#�hH�w�S;�)������1��Lm�YIs�R\�����e�e'���}�������*^�E����v6t��/g�K��R�xm�g"�l�\m��y���l�^�l�ݭ�C��g\z0$�y��C�עU������ʖ���o7�(c�����.z�vZ2����ca��ئ�
��#�?8}n,���C�����/����ȱP60��r�n�iaf�,��΋����Z@g��e�)��qML3�j{�����jd��S$����Фvv�#��)��efvI���^VgeyY��s�d�+9]������w�NT�#��L���2_-$�|����9/���"S���'��8�V�#�$����>J�H�*##�(�����ġ�%�q(G+�\����ԅ(��)j��PŖ9Yc��m��M��kq�n#���)t�kkN����]J��V=u*�O������nq���?���8|^Z�Y}P�r)@���kJVe��7�����|R?Ǣ�z/�C}��o���G��ȥ���"�^=�E"�Ȥ_��������%���~���ja�<��X���J2G[�̔eO[�#���[�B�[�ŗ�����"H;��V.JE;>���k��!f�v]��jư`��Ƞ��+��z��7s�h��`���w>�z�v��zU�Z���ʹ�d�R����r#(�FQ�D���;8D��U|�1*�J�1,��>�`���g�H��_�p�8D�&�H��E�r/��B$�)<
E	|���RxUT�rx�@��c���NO	;*N�)<$�o��N�I�c��}��4�n�u�7��t>�AsAsAsAsD�"n�g�s>�}����3�g�Ϲ�s �ND�N'��<��|e��8�q��y����7�o����4��o��	��������4�4_�4��yƄ�|&��4_�4������4�sN4��g��>6y�*I�ROV��[�loׯ��|���_=z����^Nד���y3^Lד5��y3^Lד3�ۘxuq������r�U�ȗ�����jَ!��!�������cV��&n�R���,\�͹���f��o�eHVB!�8�|�W²��T�J�	R�*P%J�m׻׻Nܣ[�[�[�NܣNܣ(p���9�m��U�.U;���/[ܾP۵)rc��q���D+D��VA�exp�[��V��K����G%r��ۜ�rI\LF��w+�w%r�(\��v�[��.)|]�K�_%�/%m��rU�v��r�7s���y/�o�c���[�xhy[U-e�iq��h���u4v�˴�ꗝR�^uԠ��-8>Zd?L���2�[$�{$���V��+/l��ǲ��y\t<�;fW��J��d�m�(�C����:��m�hf�=�����g|ǳ�c�hH��=���i�"�߱L�ئ�
���gba�h�vZ2����!���ʾ粯��I�6�����i'��I�6Rj��E��������g*���\mnG[�����;��F�џ��g���]�����)�Ϯ;�>휋����~Y�/���K3�Oq���l�!��;;c\|�$�_��ʯ�oeX��J���mv2ov�U �FA�V0~U%q��b�)7N!t���P��O���M:�rqfl�@���{���E�k:G��<*-�5�c����?�|}�3�k4�;i)�h��ФvvS�2�oʆs�d�+3�nq��<�I�t����g:����5ƚ���yYʕ�v�I���O9�J?�*#����ΦS����B�a�B�52�q�賍�F�#��^��k%y/�������Qc+�|�E�k;��"Z�H2���d�1r��$��
���<j�syN�o)���6�����_%����
I�d��>ރ��bP�P�>p����ëJ���J<��E�C���8җK��{�lR��U�6<�-���~�1�^M���M��rW�k��#�����6�JK��}X��kY��0��l%n�)v1}������j<�D��/m�N��7��-�6䝻^ۓ����7囶D�8���cVNՓ���Y;V��*K��o҄��G�}"UH�R%T��bU<�T�PS������`B0!�8D��M�&��A$PK8+�௓B$Љ4"M�yK<��Rx�'�I�Rx�'�I�RxUUUU}���'_q:��K�e�2�p��F\#.�˄e�2�p��F\#.�.h-��8-���3�d&7�Ϲ�s>�}����3�g�����O�i��?���4�柜o8�q��y����7�o8�q��y����7�����4���\.��q��u����7\n��q�-.-.-9�s��q�q�q�q��<���ƴ�'�I=*I��߫c~�|���_=z����^�z�v���&kɚ�f���&kɚ�f���`Ֆ70.��KܥUnR��)U]��~)~�\?���5�~iK�ʮ�H��w��&qKR��Lۑ9,��ۑ90����*B���+!
�P%J�@�(�T�J��[ặ�7nӷ(ӷ(ӷ(�7n�7n��/����~f�Cz顽d�V�_�6�|��jR��%v��D9塽s����_�+~_+Ç+Ç�kS
ͬ�h�P1򡹱|W�[td��|�%YB�vR�Jۣ�䫕䫈ᣈߗ���丯�q_�ۿM�GS�WS�W-�GY�wi�G[�G����ߨ��H�Ր�v�2V�f#4{M�������N��K:��P�2�C�|��eP�B�C��v! ʣ�R=��l��ǲ���[V�FkfW��J��IW̔�%C����|��m�hf�٦��g|ǳ�c��1����=���i�#�hHZ
���gba�h�vZ2����ca���*�粯���{*�����i'��I�6�z��ER�H��8>�Η�����[]������os����wwK����z3Ꮦ�q�Ү>Z[�nq�Ȓ�}Y/�Ց��Uq�����Vs�ҕ��6�E#���_�#���;'ż���6�1���l�=��T1���oeU��J��j�v6~휊ʱ�l����ۃ��|���9\e|o�PR[�x�l-��:�=
z"�����#��)/��I|�#���S�+�)��ao���x�3��a�c�I�m"���<ƅ#��g���<Ͽ�lb�[��:�^Vr��?;d�t���+B������C2;���T�+3�,W+�2T/�VW�s�/�V�������W(��%�1(pv��Gye�W���(G=�s�!DR���R��-mi�J��,�>/�C}t��N[�h=�=n�S�0y�K����ޟ���}[\_��%z�r�� ��e���� �V!#�P�[��b��:C�|�X�?~��|���<{Y_��Ի��.�|1���e9*<�f�!Gc���|ñ;�y
6J�U�D."e7Vq�!m�S����ݠj��X-�R���nȝ�����r�]�rY��M�c�Lד���U�yd���[�$��]�g�ՄiF�T�U"UH��`İ~�~�PS��������`B%P�8D��M�&��}H��($���௓B$Љ4"Y�,�yI�RxUUUUUUUUUUUU}���'_q;��\#.�˄e�2�p��F\#.�˄e�2�p��Ah���h��Ϲ�s!1�1��}����3�g�Ϲ�s?������O�i��?���4��y����7�o8�q��y����7�o8�q��y����Ӯ\.��q��u����7\n��q�-.-.-9�s��q�q�q�q��<���F�"6y�3ϱ�}���/կ��_wVO=Y<�d�Փ�VO=Y;^Lד5��y3^Lד5��y3"��`ϯvH�ŃGo"^�*�ŃGnUw�"������}]�Uە�rL�Y��M�3rLۑ9,�����nDۑ9,ܖm��R��R��R��R��R��R���������C=@�E�/��ݏ�ݏ�ݶ���ۺ��]�������[�l��d��[�n�K�֚!�-떆���f�9%�\�d��}7�<�CG*/�cX�ݦ���`�-�v]��n�C��/n�.䒮S��߈�e�ڝ��ݶwm��ʅK�j�j�h�8h�8h�{j�aR���o��*\�~�&��F�f�Sy�q~k�WXv[7�[�[�;/s�Q��n��a�k�R�C������������_�݊b*�4֢��qLF8#Dq ���ezǤ�1�+�S+�)�����b!#��1��Z
���e��h(Z
���gb`ؘ~�6����.z����穱��X|k,.{*��ʾ�ʖ|l��)5Ki"�m$U-������0){��U���q����~�{���j��Z�ǣV�j��Z������\l5돖�+�ו����Q���5�]�������Ofq���op%fòVl;3�O#rH�n�q#m����Ɋ��=��)/��՞I���|��vO�y���z%T������Ե��D%@�\�8�[N�4����4���n�S������A��!����Bځ��<LY�$��Def�#�l��c��ط����E�oal,�i���S�����,��i�v]����$���$���6r�q���g*W������P��v�6RL�������#��c��3#�Qc�eb?�����H�i�2\�B�r�����k��y!Dd|����}_~�.�B��T�+1׻��HQ%~�	/���C�,S�Ю1>4�\�-�ω�R��Ƨ�\j`ߌ_Gl���:u@��dtw�)N��k�v�o�n�#U��x1L�±�%��o��B�k!V��޿+/�T757�@�E��JlL��/ҞK�T��Z��~Y�0����Lܖ7��7�`�r�_�'j�;$��I�ܤW�Y�dSݓ_�,�VO=*��{�Y=y;���b܍qD�>����Y��Ī%*�J�X?X?X?X?X?X����8D��Y�&�I�hD���_g"�97�ɿ�M�r�)g��'���v0+�U�U�U�U�U�U'5'5'5'5'5'5'5'4e�2�p��F\#.�˄e�2�p��F\#.�˄��h������	�	�	��3�g�Ϲ�s>�}����ͩ��?6����ڟ�S�j~mOͩ��?6����ڟ�S�j}mO����>�����ڟ[S�j}mO����;�+�+�.r�r���ڟ[S�j}mO����>��q�q�q��]�]�]����������U�F2#g�<�F}���g�c=y=y=ye�������/ז_�,�^Y=y3^Lד5��y3^Lד3�ҫ#JN�����ko"_s�囋{r���y2(�ʮ��N�f�Y�Vn)�Dۑ9,�87����f��o�8pg�*��U|C"�C"�*U|*U|*U|*U}U}U}U}T�d"J��8�e�~������?؏�+�v��ۊ��+�+�{�k{�d+���D+F�!�J��(rK�[tr\�r�8s����m����{[����P2�C�J!�%
��;p���8g���"���9\-�ke���_����[tl(�;n�������8h�{j�?%��{�nn�_F���c
ó�Z��tj+�8���6h�wD?S���s�s�k.*\���~�KSj���c������l0��v[4;;�����C�0�7�~��?	 �BC��a�o��7�~v
���ja.|�۟*6�ʍ��n|�۟*6笤��)>9V?��e�K�_R�W��Rx>�O�I�6�������T��*��E����6p}���g*���\mnF�{����{��PǣV�j���ò���W���ݑ�����r����+1;�;'�#�|R;'�#�|Yč��e.P�H䕙}YY���5�go�ܱ]��s���+<�-�+2{~)#v�����ݑ�.:�
�u�:Fے�>����S8�{+	���+[~V�$��J����[�C�rO�������z,�;[�����ը[��"�#J2�c�5��Y�:dX��[��:G/$t�)�z:gE��#�_���gb9��#��>�4FG�:(Y��M�9�pa��{k(pw�+&+��I|�F��Jr_SХ������{k(G?X�F��P�JɊ�<�-�2���%$��L�+3�LW+$���݋�qY*Q�d��1��{�.��pd~��d�66��S�z�f��s���:K֮W>�sZ��h5�YQ�~��t��f�r����;Ll+��+���IT��#��Oe�vס�*ƒ۞�v,�ui�tb��{�e������Sw��d]���J����n���f�v�;l��g>
<8nR+���ձ����䚎���'d�z���k��X_�cwJ��z��׻+۶-���Ks�	�ȌJ�R���%�������	<�F#g��Y�H������4"M�B$_g"�97��<��R�)<
O���O;�
ǪǪǪǪǪǪ����������������'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�D��}���	�	�	�	��3�g�Ϲ�s>�}���~mOͩ��?6����ڟ�S�jp8P8P8P8P8P8P8P8WWWWWWWW]mO���a\a\as�s�s�\a\a\a\a\a\a\a\a\a\a\as�s�s�h��U�]�]�]�]���`F0cg�<�ʬg*�����������������)e�R������'�,���z����'�,���z����'�b�R4��Xw���dZ����"nY��'Ł;��,��'Ł;���f�8�M���Ã����J��*��"�+>�+>�CJ�CJ�*U|*U|*U|*U|*U|*U}U}T�d"J��8��؏�"��n����;�v��cum�V7U�շVv�Y�;�+�����C�^B�Q����[we-�2V��W�#�֚�͕��������&"/�J�Z�B��aTvT
;ݜ6��/Wg���]�D.�a����;N��o�o�S�=g��:��;8n�l_��/�c@ͬ�Z�B�m!���:d���!c��uܖ��#�- �����l������O;]���Ǯ�eΗ���f������k:Ե�`��0}L$-����R���j~��1�}LgƲ
�ʉ�r�j\����ƥ���l�*[+
��¥���l�*[+>�OK�K){Ie/i,��d�]��k���l� �8>�Η�����){<��k��mvr���?y���wu�Gg����n����۹\l8�~^�#��)��I}Fܗ�m�}Gs��b�6����H�)Y�g6�$p����YO���[�3�Gd�|z��,���K�$p�GZ�p4�VsY��k;|u>�I	YY����;����m�q;�tv����_)ŊS���|^�e�o��%e�!\Vw�=�^�����_�W���x�n?��i�(>w��l(],���i��go��b�7<��%@t�O�k����1W[��Ds9��d*S�;���g;FG򬒳i��{��/���h���Dd~�Q�4ҍq��I}LFG�>w9
I���Mԥ���t�y)F��{ �s��I}OO����n���J�LFVjl���O�r��q���VF��e�Oۀl��M�#���Cͺ�El���%LF��m�$IQ�D�ݏ��~K�k���#��w����W��_�&S��4*�@�_Ͼ��}Jq��5�*�~*=�K���I�&nH��Twe�)!�/
ϫ�*��g>�9¬�@������_�"��"��,��c~�%��{%�u��y�Lׯ����*K��h���Jť`ϱjش�ZQ��&|>	��D�~�~�a'����g�vp�8E�"E�"��I���R��g���M�ro�����R�)g���3���O:����K�%�Ip��R\)9�9�9�9�9�I��Nw�s�������8���8���8���8���8���8���8���8����O�i�������7�o8�q��y���ͩ��?6����ڟ�S�j~mN







��o��}��0�q���7�a���o��9y�9y��Uq���7�a���o��}��0�q���7�9y��U��EW9y�9y󗝜K1���`��6x4�F���������������)e�R������'�,���z����'�,���z���I�Փ��U��5�Xx�*�`�ܳ�r͹fݑ7dM�6�r�r�qH��f䙷"rY��'Ã$�{��ʯ�Ȼ
ϣҫҫҫ
�_
�_
�_
�_
�_
�_@�_@�!Y�������/�������A�Mۣ[�_X�V7V��]�V5���?��v,�Wd+�/�n��+�+�|W�����_(\��s��禋�i��s�����kM���K���y
/!@�d��c�!/�����ʅK�(v1	}��Wm�Om�Om�g�]g�\��]dC�/�cѱ����y�i�r�XOE��W/�#V�I]�B⻒���`a��+��
�����mv0�m�����/e��y��<�v���O�m��6���i��F�vQ�m�oec��X�v4�]�&�cI�����u���}/c'��d���������2z^�O��ȸ�9g"�kl���=��ݽ�{���6�U��ʸ��V󻑼��o;����z5a�F���\{w+�n��qb�{�+��b���/����I/�䕙=�Y�ߕ�=�Y���d��RFߑ�>,R�r�i��,vP-�
�n��d��@�v�4;>��e�Z��ⵎ>�N��;.+Y��r��F�"�-�::.�b<��V�%.��e���C�x2:;�%���b=!zxڞ�*_i�v��܀o{#�=Xww��M�R��x�J�����=�D���aeP�%�l75w;,��Q�f����̤+��pDB�b�����Y$v����%����KUƲ9�줜�[��.�ݕ�v΅%�QW-��2Ҿq�����I��R�/\���
�����oK���ȳ��%{ޑ�h�)��H�5s ���輭�V�}�#Ǡ����M;vJ�L���؋�B�e��U��n��w]6�nA�I[l�������uV]t~T�k��.����V5�ӻ%��7>^��V��V�F��F!�v/�F�G�!r�mٮR'%��U~܉r�\�h�`]�H�ۓO�X�O�M|*Ml��5ݹe����ȍ����������,j��V,���Dߑ~DM����Dk5���`}`}��
y�S�����$�?��������7�ɿ�Y�,���������I���R��g������&�9g���O9<��3���ꤸR\).�
K�%���7B7B7D�tN7D�tN7D�tN'D�tN'D�tN'D�tN'D�tN'D�tN'D�tN'D�tN'D�O�i��?8�q��@�@�@�y����7�o8�q��@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�\a���o��}��0�q���7�a������^|�碫EV���7�a���o��}��0�q��r��/>r��U��EVj,�Z*�Uh��U&�I�(Ԋ5"�Y�N��gbϓUϓUϓUϓUϓ]ϓ]ϓ]Փ]זO^Y=yd��זO^Y=yd��Փ��Փ��,����g~�����&vI��gd��"qH��f챻,nI�R'%�w,����O�}���2.�d]�J��J��J��J��J��J��J��d"���8�e�}�_u�C{�ŷuX�S��X�[wV��]MܫN�X�V;��^+����ă�9�x�+�|W�+�����|��<�B�L6�*?/����P.�"�h��n�7�v��g[��e�$��Zo��h�����iѲ���Cq��T\�n�^֧��ҁ�{X������{ky��yy��݋��G��+�t�56�H�n+R:�J���C���k! �H�6�y���k`��߿���ַ��g\kc+�lg�[c���������C��������wl!�쟍��q��n6�M��ɸ��7[&�l�\m��y���op=��v���C܈c����g����F����i{�Z�Ƿ^����xc����~����ÊG��X��o�m�|O&s���r{��O~VVxeeg�VVxqI���|z|C8�p��M�����G�J�x2�^Hq:;�����,����c�=��y���c�<+�Yjy�H~��T�u�gn���d�Vqn���Zns$B�.��#V�k�k~�Y��p�=��n$���Sa>T�/l��AHZ�S*�S"����!�e��촸�5c��F��%�������,��nB��+��W�J�/�%�;�:�r��C����
͒God����fV|oF��r�(u69%�R�������s����n��J�\=�����N��t�$���jVl�p�o����f����G��c�(�~Z2�ʯ�2P��ܶ�i���U�m�TY-�*�Jߗ����]���Kn�/�����.+컪ުۤ�j���ȑ})��.R��Eؿe���X���#*Ew�Y?����b�J���J�8�4+!ϟn�Ã~���,j���wz�`�mط�ܒyܤ��X�*�YĬ�n��ߟ'iIڶ-(�|��ߑ	<��&%"�I���I��'�|���0��������ݳ�vM���?���o���������������������NO	:�7�@��v3��걸�'5%�Ip��RsRsRsRsF�n���n���n���n��f}����3�g�Ϲ�s>�}����3�g�Ϲ�s?柜o8�q�m m m:�y����7�o8�q��@�@�@�@�@�@�@�@�u�u�u�u�u�u�u�u�s��9y�9y�9y�9y�a������^z*�Uh��U�^y��^y��^y��^y��^y��^x��Z��Ej�EV��Z*��3���O9de����ѷdԓ�RNU,��K%�R�yT�^U&�*�U�I��ɪ�I��&���zRi�I��&���zRiʫ��Ɣ���%,�`R4�������w�E=y3^XՓ��yc�Lז7e��;vXܓ8�K��vXܑ7$N+5�����p�϶U|*U|*U|*U|*U|*U|*U|+!�P4�վ?�F?�v?�v/�|7^�(�z/��n)�WӸ�X�[u�$�7��7vr�+�+�)��R�)����.Wr\�d��|�m\��\�M
e��D'��1��*�v�/��K�b�0�ژnm5FZ/qʶ�����i�w�޺�w]�cF�ۛcmͳ�c��1�b���vmE����q����[p�a�vpڸ�/ ���?u���o����[����:vi"ˢC���t�`��>��k���=��lg����H��f+ݤ�{����¸��W���[_\wd��vO#��W�'�}y���6�{"�od[��y��o7�-��y���op!��1���;�?�D���~����#��Ն6�ǷW����l5�[��/�\e�^���a�\l8�~^��6�Fܗ��H�O$����z�l����z�ns#~g27��B�fR��c�)����$�'���"=*��Kt�Y-��e�/���U+m�t1�ܐ�0��D?џ%㰭ga���e��mƢ������6�5�:�ġ��r5�	|�c[ͦ�ҁk{X���|졷*]�6e�l%�Wf��[Gʝ��l-�m*�
�%`S$��*QM��-�W� �|{aQ]L�ݓ���7h<�d����bw8��+�������X6ߧ�2D��p�~R���;�������w����ݿ;P-��o+=��We ���jR��VuemK �ɵ�n�5��]�o���d*�g�7#M�wiͩ�Z�wR��K�!Λ�W~�%p��p���Ք.Td+�oe���S�j���3ߑ7�)}+��^�/�`�R;e��ʨ�eTb3�`;dNI3�N�oȝ���Ge�J��^ՓϲO~�|�,T������_=��T��ĤPIe�7�X2,Y�TK#��U���g�"��B$�R�<"���?��?n��_�	~%�~n���&�FYvO�|��7����ʓʓʓ��������ʿ�����O��� ga;��X�N����7B7�7B7B7B7B7B'�7D�tN7D�tN'D�tN'D�tO�g�Ϲ�s>�}����3�g�Ϲ�s>�}����3�7�o8�q�m m:�u������������������.�.�.�.�.�.�.�.�/>r��/>r��/>r��/>r��9y�9y��U��5iy旞iy旞iy旞iy旞iy旞:�uX�QZ��E��EV��Q?ѐ�����e�2��y=%Z��:��e^r,�,���d�%R.rk1�Yts��*�0e�;N��J����å"��_|�5'�K#*F��,��Ȩ���׳��"���w���UWs{�3���Łw�����)�ȧr���{�m�6��f�O�U>+6��!
Ҿ�|+J�܇�ȻҫmգmգϾ/�}�^�;v�_Ju�۰�$7U ���я�+{��W*2����/(m�P۞W��W����G�~/�셹}�vv]��wR����J�I\,�k;�-���J�d��-�Z/���%m��=���?�[X��q�iַ��}D�q������m�q2Zd������m|���+m�2R�����#��Q}�u�^������ֲQ�9�f�q#H=i�X�;�2��C��E2��D���I�L�Yȑ�	<�����l�G�k��(��H�슸��󟔊G{d�ǶO��p]���g\z0+�Fq����,���|�d��J��q��u�_?�ݳ�=_/�#����僵���܌泻%�;����sY�b���c/���b�?Ɋ��ed�@�{x�
���R�~�s��}�xVs$S�
�"�����R.>��kwv;��<Wd�]�S����۱*|�,�C*��J�%K+�}c�N��ܿ[m�ߗ����[tr\�d�2WCnr�J�ex�m����n�n�n�n�*�*�"u��\��=d+6��-��g@��~Ar�a6����^�[m��Cbu?�����N�/���l�ԝ��gN��C��q>�'a ��i�����l���	ݧBG��${�w;&�G��>Z�:+[�(t�̡�[����T�ڋ/ZV��!@��ѻ�6��//����c�u�y}�6��WY
�-
�S�w;�wM�~���7�7ܮ�ܮ��+n��r�!nN��9�N՜��V��F��v/�8l�@�P0T	U�C�������O�E~��{������/ߖ_�&���{�i�ɧ�^�m׸��U�*��W�v�zV,��RO>5�ՍiF4�YX0L��������������`Y�0?�����p�8E�"M�ro��&�vM�rn��u�����g&�9<��3���O9<� ga;�@����v3����� ga;�u���v7���'5'5';�tN7D�tN'�'D�tN'D�tN'D�N3�dg�Ϲ�s>�}���sO�i��?���4������pZ/��v'�؞wby݂����j}mO����>�����ڟ[S�¸¸¸¸¸¸¸��.�.�.�.�.�.�.�.�U��EV��Z*�Uh��.ͅ�6l,�Y��ac�c�c�c�c�c�c�c�f�ͅ�^y��^y��^y��j��ի�WV��]Z��u��EV��P�PP��+�cj�RK�RK��դ��"�h�K4K+����K4`���I�RANM^��2,��ʥ�eR�tp%��XO>��MV���5'�I�x��#ZRl:�ʺRz:R��d�u���Y�����,n��r�U����*��gG�Y=+��;�$Sד5e�y3�Lݑ.X7�ʮ��Յk�µ��t���_Ã���|6UF!*����t	U�+�����(�2�*��c��^tݺ2���J2��[-� �1|��[s�Wi��k�jΛ�v��v�r�A�b�҇"RߞK�����]��I�\��vђ�'��������*�k{N번K�"�{��=��]mb�'��eͭ���ӭwm����~�n��7+����ֶq��������+m�^��aN����l��q|{
t���F��֥(��.') �I�����Q1M4/ea������W�'���9/�b����/�%��Q��br3�l�Gz,8F��J�~�"K�2$��"Gl3�L�����2z��Sr���������8�d��+2z��g�9���6�����F�+�Օ�6���W~�/��Iy�����+T	Y��e��e2��rIzd����67(b�m��2!�������t���I]�����^���:Jܗ��#=�ݔC�+��M��bv���f�#o7Vy]�����wgNݜ�r��ᗔ�-b�e�|�e�丯����r]�o��p��p��p��p�����~U�D0��Qz�Vmgm�΁��Fr�`�1ݜ^�[��CcrШ-LB'S��E�50��Ub�cM��V)4�Md7��?�e��E����W��+Φ�	��F�r𨯢坅h�\���rr�$���졸�F�/kM�~�!W� ��bvu���*��ò���Cp�(���\�*�w��w��7m���7��o߈仒۞Knr����-��wg �+z��u��t���(�po�`N!f�`!X�g8U����φDߓO�X�ϒO>I<�$��ϒO>I<�$�ܰnX7,���,o챿���*I�RO>6y�ύ�Dc"1����������������$��p�8E�"�g��;?��;?��;?��v���?7l�ݓu�����g&�97Yɺ�O9<���������z�z�z�z�z�z�z�z�z�z�n'cq;���N��t�Ԝ��|n���N���N���N�����h��Ϲ�s>�����C������sO�i��?���4������pZ/��v'��-��?���q�q�q�q�q�q�q�q�q�q�q�q�q�q�q��]�]�]�]�]�]�]�]��EV��Z*�Uh��U�6l,�Y��af�ͅ�]�]�]�]�]�]�]�]�6iy旞iy旞iy旝��WV��]Z��uj����Q���Z*��! Q0�c`���a������V6
�$L�lX�*�{�2/2)=ńe�H$����/���s_���6����g'�g'�g_/"��&��'���
vR�	|�6p,'�_|�O=)e��+�U�)4�%R�zX���q`K�W�cRz9��r,/��`ذ),��^,
���<��;x2�Vtwd����r����°j��Q���?��2.�t��5���.R$7V�7v�7V����c����/e۫[�;qM�_N�Cs���x�{�D�`)��d-�r�;vt�ġ�vJ����%�.K�w$��|��G;�)r_�ᣈᣈᣴ���Ӡt�7s��v6�[���//�n;��z�m��7��/�M�w{������҇d���O�*�'�����Y`������9^$���S��$���N�� �d��2%jB�O����/4*&���kdد�Vj3�ug�9�k��rj^�E#��^<�r��	T�����MY�Ւ�}\�a�#�\__�����7��pK���qIz���qq�����d�ef_W��qgM�)r�2�.)�#�m��ߑ�M�:��e��yn��۩�^F�B���Kr����ܶ�+M�]�n�v�j+v��/))`Sr+wg��Ȝ��l�!vU��*Ӳ�S��b����vQ��RA׾A׾?���"�J�����9/�җn<��Cv���]�8�K�m�:m�:n�����oߝ᫬�Z�D4l��Q��*g@��B�6��͝�[m���l61zMLB'Y@��E�5��̴6Y��S�u���D+�Z!��@��C~�h��W�7�D+����+�q���r��8��yo�x�9]��0�}�Fw���/�-�WYí�\e�*졸��:ȆdC�!�S
�����oߕ�#~�F��^I�y'%rO%�<���W+���/ueݝ�vv]��{.�{.�{.Ӵ���(�po�Y�,ݲ'l��"p��f��|2+����6��z�`�X.V���b�X�,���^�z��פ��$��'�I<�����>6y�ȌdF%PS�AO����x0����$��p�8E�"�g��;?�yH��P7Ƞo�@�"��E|��7Yɺ�M�rn��u�����3��ο���ǪǪǪǪǪǪǪǪǪǪǪǪ��v7������9�9�9��q�'�q:'�q:'�q:'�pZ'�s>�}����C�����ИИИИИИИИ�sNE�<��������
�
�
�
�
�
�
���������������������Ϝ���Ϝ���Ϝ����EV��Z*�Uh��U��6l,�Y��af�ͅ���������6l,���/<���/<���/;WV��]Z��uj����]c�<uX��u��p����K��R�h��Q������_�����gcjM_ξ�4#cYWVU�_#�~9�Y<m��7�#hȬe��0ȩ0��h��N2,��,��&���&rhĊ5�a<��V3�I��ɥ�$X{$Xt��s�/��`RQ�Fݓ��a�c����W�`������aG>��E��Ԋ	"��I��Y�������ɁWnΎ�^܌<9{s��I�V-���t���Q�qh�na���y3V8��x��\���n�3��ʼ6m�Eʽҫ[�c�na�iN��}�~^J����q�w*�;�ʲ����j�b��v��vP۵ʶ���"r\��-��(�1Z��m:gX��G����{���V��_�ҁ��'Sr��o+�����\kc�^�7�N��oڦ��v��� �z+�q��l_�ʷ���d��v޵�l%>��[���2�dcg��i[2��8�8�7��+$m��Ց՞Ζ��+1=���#����_W��������Vw%f'rGe8���UKg&�)��,w�8��p���'��V{8�#�ǭv�NNH��i�W'���u�V�
�����vZ�'��ܕ@��=��&����P+�\���F����"A엏ʑ	�f�jѦ���]��#���:ܩeҾ��|^�)qZ��"�7�V;]����8��8������[��\Tr�tq�q�q�q��v��r]�v����ۍ�_��/�g��B�v1݌B7[����vq��^�e@��Ccv��T^';@����l����fW�β�c���#v���d6Y����yV�ݍb�im���"{�g��ʠs�o��0�i�vv�z����?�gm罧u�Cq��0�}L*_S
��~U�pݒ�җP�I[i*�<�%Ĕ8��������s��%oI[�SugM՜��v��v/*���!f��8d��c�X�9+��w$��,rK*��rŹHܤnR7)����e#���H�jƵcZ��X֬kV5�<��Dc"1*�J�R�)��`B0!�F�����E�"��H��_�/)��&�I��M�rn��u�����g,�K.˄��,�K.�U�U�U�V=V=V=V=V=V=V=V=V=V=V=V=V7������9�9�9�tN7D�tN32222223�g�Ϲ�s>�}����C���LhLhLhLhLhLhLhLhLo����-�h�E�sO�4�������9w9w9w9w9w9w9w9v��Z*�Uh��U��EV��Z*�Uh��U��EVl,�Y��af�ͅ�69v9v9v9v9v9v9v9v9v9v:�uX��c��Uj��ի�WV��]Z�}���<uX��s������o��/���?|�����n���V�'����P^Q�V�k�h��Ѱ��cv'��
��ڲ�2x�V0Ub|�
�c	v���?ѾV0���$�&x6dV7��NE�D�E~e8ʶ0�i?�|d
'�'�2��'�VOvYFYvMv����6�IW����_vO/�_G^����������FKvE=�U]�UX��8�:o'Z���s_r�cnշ��7_CJ_�N��҉o�݆�ڠj��_ۀ��ѧnf���¥W�٢3��ы���?,�܉ӵp�!_�0��/:v��&9K���/��u�B�i�]vu���ceݗ���1{�7~�Rw*�a���[ȣ �Q�qs���v���n�$N�c�qʶ���bu����l�B��ӡ6��(��M;�����H�~��pT��%Xbm�2����HrU|Si�s���}�Y#m�̞�)Y�p=�'r�;|vN���.Y�'�Vj8��f�{;a-�^s�M˥�P8	��P<zf�#qt��U@�D1I��"����H��}o8�V�n�����u�����+��������c�p�1{�"�2w%�~��"Cr.�5���q�5��s��3��y�s���H��P�c��-����[ug[ݣMܫN�N՜��~/�r���+�ܕ�앷G%r��ۜ��G�/���h�P:�!�;l&�����e���Fl���f�!��Fl��**/���ga_�4�Kln�?��y�P �1x͍b�im���cu0��d^�eX���k�R�/(K7�؝d+�w��w�#��!kY@Ǧ��Z�P1�%�ݵe+��G�G�G+�w%�9C�e�H:�^����.ąؐ���u7Vv�R�*V%H��m�[r�����po�`_�"p��w%{���^�\��*�ܝ�`ݱvR5�Z�xּk^5�׍k�5�Q�(ƔKJ%�҉dF2#��Ī
r�)ʠ�����������������������"��K?����)g���Y�_�_�_�_�_�_�_�_�,����rˉ�.'_q:����N��v�ԜԜԜԜԜԜї˄e�2�p��F\#.�˄g;�tN'D� � � � � � � � �>�}̄ƄƄƄ���3�g��LhLhLhLhLhLhLhLhLhLo����-��8Lo8�e�������������������������������*�Uh��U��EV��Z*�Uh��U��EV��Y��af�ͅ�6l,�X����������������������c��U��U��WV��]Z��uj���ߎ��ў:3�Fy���@��������%���@��y�������y��E���� y��u�����&�/�~�>��7��){��_������ۋ��_��p����Fѓ��I��p��I�ݓ��	�p�/��~q��Ђ�8�w���������y?�{7cz�'���Y�"�9��!�D���%�HȰ�Y�'�g��"��&�ɑ��������nUwnUvَ�ց�qr��ϤI��_�V.)[�]�;��]��)5��v�"U҉k�7,Q��E�X�]�n�H[a���e�n���V^/�F��j��V�����P"c���:<�m��oW�;J�r	�߱Cp*�0*�W�#[��V��i[�����|��/%K9Qxv{�M���Rm��^W%��66�e����1u�T*�����r��(�JOl�dTr�(c廊��Y�O���B��@�i���#�<2:F���VڎV�F���r{�|VA�d��G��2�_ǭv�~Kv�S)�#����w�Û9�V �-���m�,�D~�QN�l#�zĊv�1�{d����'CeTaR+�2'$�r�m��2$BU/m��m�]�i]��ն�N!'P,սZ0�;J��|�������ug�P0�%�Jr���������7'(nO%r�%m��o��xq�4k?:�?:�? s�p:��M�������Y�	���B����NTC�v����Bm-���n�������"u1�G��G���B'S��Ӥ��,�/��r���-[���ܘe�W��Z�R�-
é�f�m��/ �.+�+�R�R�%��[�UM�Yu�]T���s�z���d)�n
/������N/�8���`_
��l��'rW�+ܖ�{���`�W�V�틲��Ռj�5c��XƬKV%�ωgĳ���L�&|U�D�Q)TJU<��F#��������������g��I���R)<
O����*����������������e���\NYq:����N��u���������挸F\#.�˄e�2�p��F\"tN'D� � � �>�}�����7�hLhLhLhLhLhLo9�s<�y��i�����O���?���i	��4�_����	�i�]�]�]�]�]�]�]�]��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U�6l,�Y��af�ͅ�]�]�]�]�]�]�]�]�]�]��V:�uX��Z��uj��ի�WV��j�����<tg��<s���t`n.��v�D��U�֍�k�cu�w�[��պ���q��ӝ��n��:y����4~�������i�Ɓ�����B��Td
'��4&�&d&d����s�s�s�\a@��;�Wa4_��؞�c e� j���������Ip��FsFsRuXyX�K ��+)U}�=\���x�4\�1��/��`Ʒ,����vu��ʣo)?T��UҰ�V��%���Y�$�R����E��Ҍ`�n�]ߑf챿#��'��O>�G{r�r��?�qm���g/���`ui}n�Q܍��Ճ̓Ղkĳ��>�c���U�.���	���l��8����T~�g[�JW+�^_�[��H5�ؼL�)`�|�D�PJ�E��m:Ɵ���S�d<��SSg���J̟o$Cx�"�HЬW'�+$��A�"�ig��G�!Pb���r|>=*��ҭ��go��G�
��Gk�e�ov�W�9\]-�C�����v��nP�������^�;�2y�K2y�K2k�2+�X�2+�VzF�cr��&�
���,E�Wk���dBL�Y�R$CϾ*P0P�R?�|_=�D$Kn
�*H9��NBվB�HZ�]!k�}���.�%�,2W�+�ԕ��J�ѝ����p�b9 r�}q�9n�L�o�O���#��S��[m��Ӭ6q��J�q���߄�o�d�����{~�P[:ܳS��[cr��^˶]��v��-t��wS
͋잦����\��sYu�]U�]!k�.ą���%7=N�S����bT�J��R/����(��h���R'��,v�:0���4�%��z�^�X.V+�r��`ܰnصiQ�X��KV%�ωg�3���L��&���������՜"�"��H��_�/)���E�"�yI�Rx�'�I�Rx�'�X\,.��5�5�5�5�5�5�5�5�5�5�5�5'5'5'5'4e�2�p��F\#.�˄e�2�p��D�N���N��fAf}��i����O��m>�BcBcBcBcBcBcy����4����������o���4�����i�]�^|���^|���^|���^z*�Uh��U��EV��Y��Qf��E��5j,�Z*�Uh��U��EV��Y��^y��^y��^y��^x��c��U��V:�uV��UZ��Ej���+TV��]Z��uj��ի�ڻ~:3�Fx����Z��iq���.��v�5��Ϯ��t]�y���	�����\��F6�Mٰ�Zc�c¸�}Ɖ��w�;��ם����}����Ϝ��7���m q��}̄��i.�U��5j-Wo��G�17�.�*�p��E�sO���(Lh-���p����p����D���e��0�#.�XaȰ��cVY��Ru`XO�Fޔ}���&�p��򳉞�\��ϳ�B$Љ�ɡ�*Ni���Uv�I�&�ω�"�X�J�X0I7���M��r�Z����&�"��ω��FM�g�	V��"����;?,�[���F����nZ��[n�=�_W�o���{�5�����D�y?�i�)CnV��^���������?���Y�}�� ���W'@���l���7�~��H���f"C��oh�d_���=��'�V>;��?)���o���{-�����������Y��+6����8k�ߓ�ߖ_�׉m�O�EG�E/��X�V�z�'�nY$����j�v?�W�N�`_�]ᓡ�7�0'�D,�_"q|��0T4~�N�Sr|�W�t�eҜ����$��Jr����V�J�.}�CVԕ��S��M��J�\J[�$��ƛΛ�w��q������z+u��m����+��M��M��%��J��v�gb�:ܚA�͋�ѝ��70�ug(vQ�t�܆Wn^���ra����x�*ܩM�H9�.�˥;.�A�S�ՉR�*V0Q|_��6��G�.�0/�Y�&��Y>�����@��
�]�_�,m��+��r�nط,�*��X7lZ��(ּc^1�ҌiD��ZQ-(��#���`B0!����8E�"E�"��H��_�/)���E�"�yI�Rx�'�I�Rx�'�X\,.��5�5�5�5�5�5�5�5�5�5�5�4n�n�n�n�O4O4O4O4O4O4O4O4O4O4O4O4N���N��fAfAf}��i����O��m>�BcBc��i�������������������o���4��@�@�h��U��EV��Z*�Uh��U��EV��Z*�Uf��E��5j,�Y��Qh��U��EV��Z*�Uf��iy旞iy旞iy旞iy��U��V:�uX��Z��Uj���+TV��QZ��uj��ի�WV��j�����<tgj�Viy��;Wta�4��K�Viy�w�j�sU�j�iy㪵Ej����TV��QZ��E�]�^z-9ڻ��a�4��ў:3�V����/;�+�+�M���uĺ��⋜��վ��(�⋝�;�w^j��Y��y�y�y���.�ii	�������\З��('��~����o�FU��]�������Y����Á/_	F��B��I:���K�e�Ip��R\).������ap��X\$��~i=�Op��%�)d
Y�yI���Ro)4
M�u�����o�u�Y��fk���e���.'&�97Yȼ��p���WԪ	��A4�'����Q�`K��/�Q��h�nȄ`kƵ���FK��e��;*�n5��F.M�¾=���������{~J=���|�}��oe���HZ�m�N�cL���#�=�d���>�)md�m+-�N�]�I�����{<�W��ۓ�ߖZݍ��I~݄��n�W��aGn�{v7nV-��#�6|T��%�+ʒ��	�X9,������,p��2�l��"vɟ�hT�
�"hm�?f�٭�n
�*V%JĩX�St���η�:vB��}7>샥F˫���B��)n��n\I\]d�.�-ˉKsFWo�Wo�Wo�Wo��r���W.,�..x��x�޲�/�̡�	(\��e�I+~%��R��e�� �Q��Λ���+y��)�W�:��:�i����η��୲���G��^��G���6��Cl�9�,����}����'�'��{���	�׹,+���^�qW��'��'�vŻbפ��kV5�ҌiF4�ZQ-(��K>
r�)��`�J���	<���;8E�"�"���Y�,�/���M�@��)4
M�rn��u�����g&�9<
O����)<��3���O;���ÚÚÚÚÚÚ�B�BÚÚ��7B'
ғ���2�p��F\#.�˄e�2�p��F\#9���,�,�,s��8,s��8,s��?��m>�}��i���7�o8�q�p�p�p�p�p�p�p�p�ڜYwYwYu�V��Z*�Uh��U��EV��Z*�Uh��U��EVk��Y��]f��u��5�k��Y��]h�=gέ��ߚ^y��^y��^y��^y�玫V:�uX��c��Uj��U�+TV��QZ��E���ў:3�uj��7�󗺗������uj�Viy��~iy旞iyڢ�/=o��F�o�/;TV��QZ��Ej���+TV���f���7�w���0ߚ^x���F�j�sU�5[�a���Z*�K�Uh����������V�uo��;�3�����u���Y��?2�2�2�2��^e��p�p�ڟ�S���O���NhNh.����3��ca.��U��v��2��a�'��'�/c��g�h�������>o��F\#9�p��|e���Ԝ���}'5���9�4_a�a�I�a�c�_�c���<���`U�V=U����;��(��,�VY��~���(��_��}��o�yH��_���?�p�8D��E��c}ʾ�e#v�r�K�I�ȿ�#�7l������P���h�qf��a��bj{Kg�]�m�����L[ ����(U�P����)��v�ؙCv�7J���3)���H2-�bO��۱qX����	W=X���j�U�å~�m�Q��R_�cwn��ʒ�(��F�r1�⍟l��gr���I}ʒ����^�o׷��2w��'p�ݲgl��&B�HT�
�"hm�?f�٭�n�*V%Jĩ[ϝ;!N�V0T�T�yi��ky�l���.��޲��ġ�q�ܸ��y�[��-�r��KsD���P�͋�ǋ�ǋ��!v\HZ�d~�^�w�/s����r��m�J/��޲�:n}Zt�u�bT�`��
�E��+��ky�J�X�-�n
?f��#�h��/"P,�	�"P$HT�
�!R$*M���d�e�����'�����'�a=�	�R8�W+���_>*��Wϊ�{�-zI�ƵcZ��(ƔcJ1�҉iD��*�����$�>����p�8D��E�g��H��_�/�7��&�I�Rh����g&�97Yɺ�O:�������������������ÚÚÚÚÚÚ�B�BÚÚ��7B'
ғ���2�p��F\#.�˄e�2�p��F\#9���,�,�,s��8,s��8,s��?��m>�}��i���7�o8�q�p�p�p�p�p�p�p�p�ڜYwYwYu�V��Z*�Uh��U��EV��Z*�Uh��U��EVk��Y��]f��u��5�k��Y��]h�=gέ��ߚ^y��^y��^y��^y�玫V:�uX��c��Uj��U�+TV��QZ��E���ў:3�uj��7�󗺗������uj��:�uY��^y��j�Viy��~�7旞:�TV��]Z�}��WV��]Z��E��4��a�����]�i�^v�ݵF�7q�ߚ�����-4Uh��U��EV��g���(�(�(�(�(�(�h�h�˼˼˼˿˿˿˼˿�@��/�S�j~q������3��'4Y�����g���e�ь�}�ЄЂ�D�F����?�Ah�l��n�y����w�����wby���g;�4]��|f�����v����.�s�7D�9�I��˅���z�z� gc��cq8޳���qvǝtk�U�͆�6L�i3Q��|nk�tNí�3���O�@��R(�a�cp�yg��J�yIW�Dc%"�ݓ�쯵_p챿M�wqz��(��z���a!gֲܙLGS;�蔵aYnRş��k�E~D
��������U���ݤj�6�uc���
���l���)TM��ڸ?ZQ.����߻~�m����FOv%�=��ܢgr���e�q���_r�����`�X�V���{n��^�φNᓻe��O�D�I��H�	2"�6E8m�/�8�
/����_�Cl�|	��.�ph�%Ud]�]�[.�[.�\^�Y��B츦�f��Z��Z���s��9�i��܉zn~�vG:�}�7K�7^�� �y�{<�[���7_�o?;��v�	����	��Q���ʮ��H���(m���٨j�@�D$Ȅ�@�!R$*D��_�&��M�����|���W߷a=��*K�T��X7l[�-����7�X߻awv��kV2z��ύ�Dc"1*�J�R�)ʠ�*�����0�������0!/��;?����Y�,�yK<��R�)g��'�W�W�I�g'���rx���'�|���x��X��z�z�z�z�z�z�9�9�9�9�9�9�9�I��ӱ�:Nw�s����'�i�q:'�q:'�q:'�pZ'�����pZ'�pZ'	�	�	�	�	�	�	�	�����3��p���Z�%��Z�%��Z�%���?6����ڝ��������[S�¸¸��.�.�.�U��EV��Z*�Uh��U��EV��Z*�Uh��U��5�k��Y��]f��u��5�k��Z(�E�:�旞iy旞iy旞iy旞iy��U��V:�uX��Z��Uj���+TV��Qc�<tg���]Z��{��|��r����+TV��Qc��/<��Ej�V:�uX�QZ��v�Wo�v�Wo�uj��ի�TX�K�F�ڻ��Zf���ڻF�����V��o�/=o�U��EV��Z*�Q��3�UqEqE֬�՟Z��V~j�̻̻̻̻��/��2�5g֬�e�ͩ��?8�q�m m<���p��8��`o���a	V6�+�&����������y�|oZ4�n�����-�h�E�Z/��|Nk�s_������'5񹯍�|nk�s_�����h����w���oY��F�F�F��oY��]���Όo:2~r��*��I��nk�s_�pY�7���UT��Y�&�uW�XyH��>6���܈�	��g>�f�Y=�l%�w���is⯞��%}��Y�l�Ү셯��`ܓQ��`ĵi}*��F�"[�{�,:�*K�lnɼ�PS����'����&�##�>	�҉kĵ�Z�M�ؖ�Kv%r���&w(���_�~�$�l[�-���r�m׶�������|2w��,�����$��$��@�!�)�l�|	��P�7@�(%L�ȧ���V��������η�q �������H:�)���������UZܪ�nUVۃ/m��m��m��X�h�g�i\S��kz�i��5�^����|x����qy2/"P$J��N/�8����5L�H�	2�"P$���"dBX�;e�c�Nᓸd�;�O>I<��'�a=�	ܬW*K�T���Ov�}���Gdkv�{��ܱ������c'�ȌdF%Q)TJU��J��*��$�a'����g��Y�����<��R�)<
O9<�Rx�'�W�W�W�X\+���������'_q:����NǪ�c�c�c�c�c�c��������q�'c�v9�I��Nw�s�7D�q��"tN'D�tN'D�tN'D�ND๠�������ND�ND�1�1�1�1�1�1�1�1���3��p����8KS��8KS��8KS��?6����ڟ�S�¸¸¸¸¸¸¸��jwWW\������*�Uh��U��EV��Z*�Uh��U��EV��Z*�]f��u��5�k��Y��]f��u��E�>uo�V�uX��c��U��V:�uX��c��U��V:�UV��QZ��Ej���,tg���ѝ��WXoa�xo���r��^�㗝��4R�Xh�Uc���Wp�a��E/u/u���+Wo�}���5���u��5�j-\��]mO���af��v�7ݵv�tn�<�o�/<���U��EV��Z*�Q��3�Fz(�E�9y�a���p��.�.�.�.�.�.�.�.�V~j��Y�����(KS��?8_�!1��AsD�#:�6�4id�J��3�����	�	i�]���'5�cz�2���-�h�E�Z/��|Nk�s_������'5񹯍�|nk�s_��Nk�s_�q�F��oY�\#.�˄e�2����w��_�����Nw�s�3��:'�I�Ip��X\$��~ie�Op��I�pWʢoύ�|l�#ZT�eT�uk���Kȿ�`�rl<86�d�򨔪�~�|�C�B۱�Cpt�/ұ��*��R_"�j�Q��I��l(ʢoύ��vM�gҤ��FE�g�K Ro,+�Q7p>�����*��|�>�>���~�W��~�v
��+�"n�D�܌�dkV5�פ��$�lW+��r�\������|2y��϶��{�%���N"B�HT��D,Щ�L��;e��d�Rk�+�	X���6U�ۑ�?�Ν�qN��X��X��m�c�ʱӥX����5�Vn��^"���������m�\[pz�2:ӳ�m�#�6�ta�+�	b,Ce����&B���,��]�H����I��5��g��gl��,v�ݲw{~��^ۓ���u���{n�{���,oݍ�v6����#ZQ�(ƬkV5�=x���o׍�"1��ANU<)�}`}`}`�Ov�g�v�"�yH���o�y�Y��<��3�������*�����������_q:����N��u����}���'Ip��R\).�
K�'5'4n�n�n�n�n���n���n���';�9�I�����	i�����3�g�Ϲ�s>�}����3�g�Ϲ��ИИИЖ�	jp��	jp����?�g���%��Z�%��Z�%��Z��S�j~mOͩ�a���o��}��0�q���7��v��o��9y�9y��Fz(�E�=g���Q��3�Fz(�E�=g���Q��3�u��5�k��Y��]f��u��5�k�g���տ�[�ў:3�Fx���<tg���ў:3�Fx���<tg���U��TV��QZ��Ej��<tgj����o��/|��z-]�/<4R�Xh���E���㗝��4R�R�Xh�Uc��k��}���5���u��5j-\��]mO�5ŧ9u���}��ں�Fx�K�4��Uh��U��EV��g���]c�<tg���o�j�[W`q��/>r�������/5g��՟�/�_�-O���HLo��\ѝg�q�7�>�Aa�����v��&���3�7�w��ItNk�n.�s�BD�_��-�h�E�9���|Nk�s_������75񹯍�|��_������e�2�p��F\#.�˄e�3��������꤁�$� gc�c���\%�Rn�gU'T�&�I����Ҥ�%�c/�cW"�^UIG"6y�(�|KJ6���U��x�9ZQ7°��cl��������"�g�Ѱ����"��M�ro�B_g|����X0Wȿ��)7��#
�W��>�E�g������
x?X�쏭(F���������_�~��Q-(ƔcV5�ݤ�#��r�\�\�K�{~��`�m|�k��'~K'�,�*D�H���L��;e��c�N��N!&�
�Q�`Z�`�ʳE�4E�4E�4G�Y������V:������n��^ہ��&��c�ȱ���E����.#���l��?��/gj!&�@�_�N,D%�T��,�*M|*M|*M|*M�}�w�����ݲwl��^�p׹,��z�^�X.V���`ܰnX7i'�I>���FO�2}��ωiF4�Q�X���OV2z���D�Q)T�~�>��p�8F����ȼ�^Rh�&�I�g'���u�U�U�T�
K�UUU����c�c�c�_q:����N��u����}���'Ip��R\).�
K�'5'4n�n�n�n�n���n���n���';�9�I�����	i�����3�g�Ϲ�s>�}����3�g�Ϲ��?���i���/�_p����?�g���%��Z�%��Z�%��Z��S�j~mOͩ�a���o��}��0�q���7��v��o��9y�9y��Fz(�E�=g���Q��3�Fz(�E�=g���Q��3�u��5�k��Y��]f��u��5�k�g���տ�[�ў:3�Fx���<tg���ў:3�Fx���<tg�����TV��QZ��Ej��<tgj����o��/|��|���j�4Xh��Ϟ:0<���~9yᢗ����E�^y�ߚ��_~k��Y��]f��E��EW9uŧ\n������|�]���:3�U���EV��Z*�(�(�(�UZ��Ej���ߢ^�<4n-U뚮iy旟9y�9y�9wYt���V~e�����i	��2D�n�g}'������U��F����Q�PZs �>�}�8+W�h���,�Lo��s>�}̂̂̂̂̂̂̌̌̌̌̌̌̌�8�s��8����'5'5%�Ip��R\)9�9�9�9�y�y�:�<����o��]��]��X�����RΩd
M�,�K<�Q7l௓�H���.ܤV�$��p�۲�J95t�n�F2 �MZJ�~��Ս���J��)1��a�AQ��W�XyAaX�3�j�:�z����������l<�.�Y5d�)?4�������Y�}H��q3���՜"���#�#�#�>
z�g�~���L�ƔKJ%�ՍvF�i'�H�m�9,\�-�	��φ�|6����϶N��O�L��!R'��&v�ݲwm|�$��$�aR*0�<=�x�X:"�q	W8���E7�7�6E�g/���Ȫ��Ub�*�	5��M��&��h�����Cpn#�<��!�,1	5����p�b!,B���=�e�T��*Yv,��'���}���m|�l6��~ŷb�qX8�V.+�vŻbݱn�O�5�=X��D��Y�L�&|J%�҉g�]ό���������g��H��_��"�yH���)4
O:��<��3�����椸X\,.��5�5&e&e�5�5�5�5���4_a��jK�%�Ip��R\)9�9�3#3#3#3#3#3#3#3#tN7D�9�I��Nw���hKH,�,�,�,Ϲ�s>�}����3�g�Ϲ�s>����i�����O�_�����p����?�g��-N��-N��-N��ڟ�S�j~mN��o��}��0�q���7�a����o��}���Ϝ����EV�3�Fz(�E�=g���Q��3�Fz(�E�=g���Q�k��}���5����ߚ��_~k��}���5��wEۼ���F���WV��]Z��uj���:3�Fx���<tg����Z��Uj���+TV��Qc�<tg���]Z��{��|���F�Ѿ}tK��G���Z�͆���|�Z�j�9yᢗ����E�^|�]�uj����]f��u��5j-\��]mO���Zs�a���ں�uj�V:�r�Z*�Uh��U���EU��4V����-Q环\r�q�旞iy旞iy�9y�s�\U@�y�?2�2����?�BcBc}̂�8γ������O7i:Ѥ�F���H��D�}̄ƌ�|Nk�_��f��<��Ɓ�}����3�dddddddfdfdfdfdfdfdfdf9�c�n���n�'5%�7B7�7B7B7B7B7B7��B������O�DݓFёRU����I���Ro)7���2������(F偎�Ñ�'2Eϰ�ϰ�հ�*�dA5lo��a�,�ό����"
�DM[��1��0-Yg;?�l.�*8���H����I�Փ�ap��Y���/,�̖\0?�P)�Yp�B$�R(%�L��g"�Y�,��F��G�|�য়9TJUȌiD����X�dkv��H�qR.V+��~�{��p�;k��_>�;�Y?�d�$�T��&v�ݲw��k�j1:��)~�<q<Ь�t<�	�BE/@�K�%�bʰ�e���*OF�&��c�I�P$١�-{>tp���8������*Yw�Y8��p�5�2y��/��]�H�¤TaR˿�{�k��_>����8l6������bݱqX�l\V-��vŻbݱvF�#Z��҉iD��YY�L�&|J%�~DM��p~�>�>��p���E�"�yH���)4
O�������挸F�F�RsX\,9�y�t)3)3)3,9�9�9�9�4_a���s�7B'�7B'�7B'�7B'�32B32B32232327D�tN������|N��Ƅ��̂̂����3�g�Ϲ�s>�}����3�g�����?���i���/�P��	jp����%��Z�%��Z�%��Z�%���?6����ڝ��0�q���7�a���o��[Wn0�q���7�9y󗞊�g���Q��3�Fz(�E�=g���Q��3�Fz(�E�<�Y��_~k��ߚ�5���}���_~k�n�>th�}��WV��]Z��uj���:3�Fx���<tg���ѝ�+TV��QZ��Ej��:3�Fx���ի�7��<7�^�Ѿto��]���q������ٰ�㞋M��֪��K�K޵u���ժ��Fx��5[�U��ժ,uX��Ϝ���Ϝ��U�5[�U��;WV��Qa����7���{�7��f��iy旞�7��~�7��\�n1�ц�uV��QZ��E΋�U�Uĺ�]��[Ho9��>� ��3����l!*��ձ��I֍$��7���e��ˋ�2�8^p��BZ��w��8-�h���h���h����D�F\"y�y��#t).7��|g;�9����w��]���qv���w�\"tN'D�>�BZBcR\,`VU��ϷȢh��U���'�K>�Y�rϳ�D��&x��F_�a/�'��'�ȱ�g��k�����"�H��q+8�bUȍ�Dl吉d"M�}����Љg��������c��RuX\,.�����'�I�{���_�_�_�'�I�{���Y�W�K?�Љ4"M�A$PI����	*�J�Y���	���`�0`�0L�&�c^1�ݤ��r��_=�	��/����'��Om|�d�;~��,�l�}����'�,����,���q	���E�"�@�c�������I�D$֢kP�fT�䲌*O/�'��I�B�Y�R,ߒl�l�l}��]��_�k_�k]��0�5_�e�5��5�e*���ϊ�|U�ۯo׸k�5�T�
��U���~X;l[�Ke#V��HդvR5cZ��X�|K>%�ҌjƵcZ��X���0~�~�~�~�>���>���>���P�ȡ/�B_"��E	|����o����rx��X�N7��9�.<�:'�s � �#3#3#3#3#3#3#3#3)9�I��Nw�s��������h�f}Ђ�����23�dg��,Ϲ�Y�s � �>�D�F��oY�hBc}����3�g�Ϲ�sO�i��?��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	����HHLo8�q���?���4�������O�i��w�k�8��|;�ڟ[Wzڻ��EV��Z(�E�=gq���7�a���o��}��0�q���7�a���o��}��0����v���G������j�<4yڻ�o�/wF�U�4��U�5[�]Z��uj��ի�WV����{�7���{�7���{�7�]Z��u���旚^iy�旚^iy��Vj�U���9��v�5�-1˱˳ah��i���V){��K�K�a��E���Y�<tgj��ի�tg���Q�:��~j��<tg���]Z��uj��<tg���ў:3�Fx��V:�uY��^y���0��5[�tta�U�+TV��Qs��Uq.��\K��u��i���2����07�y��^2223�7�o���!1�1������E.u`�ՄƄƄƄƄƄ����2C�d&4&4N4f�o5'7�o��q�� � �"tN'D�`j��դ�F��ۋ����|O5%��a�_�,�|�
�e[8ʴ�T�T�T�T�T�*H$2���U�r,n�ĥ��7՜K1���H��o�d"O�_�_��K �ϳ�}����������+++�
�ap��uK:��RΩgT��Y�'�I�{���Y�&�I�Rx�a�,��K?�Љ4"M�g������J���|l��g*�J��Ī1�ȌdF2#��X֬k^�}�7���v�w)=���p�8l�.K݋n��`�rX.U�z�^�W�U��=�����y�<��^,�
�a�K0�$֢kQ	5����*Y�,�
�a�K0¤Y�R,ЩhT�7���l���_�O/�'����������W�r���c~�������`�o�8k�5���~ſH�qF�^1�҉iF4�ZQ�(��c#�"	�ωg�4�Q-(��
r�)ʠ�*���0W��_�}�"�&�97�ɿ�M�ro������7������3���$�g�q�gqv'��<��|���';�9�I��Nw�s�������|n���';�9�I����7cn.�f}����3�g�Ϲ�s>�}����3�g�Ϲ�s>�D�F��oY�h}̄����3�g�Ϲ��O�i��?��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	��
����7�o8��O�7�o8�q��y����8��[S�j}mN��o�/>r��/>r��V�uo�V�uo��}��0�q���7�a���o��}��0�q���7�a���oц�oц�oц�oц�oц�oц����/<���U���ի�WV��]Z��uj��7���{�7���{�7�޵uj���:3�Fr�K�/4���K�/4��f�5Y�͎�F�1Ѹ�G4���c��/<���U����{����/u/u/u/u����tg��֮�]f��Fz(�E�=g���]f��u��;�(�E�=g���Q��3�Fy��]f��Fz(�E�:��ګ��{�(�5�k��Z*��s��������.�.������M���
��L(L(L(L/����2���P5P5^e�2������6�	�	�	�	�	�	���4g�o��s"q�3#t)9��"q�q�q�3#3#3#tN7D�tN7D�3#3"q�q�q�s"s#4).=V3��}�&��&��
�
�
���g,�H��5{$ٷdZ5d��,j�F_g9d"Y�B$�Ro�E�A%����4"E	|��7��<��Rx��g'���u�U�V��rx��g'���rx��g'��UUT�rx��g,�|��O����)<
E�"��Y�0>���_o�AO"&��˺Q�t�h�Dߑ~DM�7�Dߑ~�M�Q-(��d�#'�I=���.�X]�I�᯿����	��O~�w+��r�\�+���`ܰnW�,�K
<�w������d�xd�xd�xd�{e��e��e��e��e��e��e��e��R,Щo�6?�6>�f�f�f�fK
<�y+�䯿n�{v۰��^ťbױkطl\V.+݋���`ߤrX��Q�⍟dd����L�)��3য়ς�|U�B%P�T##�#�#�>
r�)ʠ�*���
r�)ʠ�*���
r/���E�"��K<��Ro�yK<��V3����� gI}$��7���oY���e�2�cqv�������7ln.��]�����q�'�t���}';�9���3�g�Ϲ�s>�}̂�8-��8-��8-��8-����q�g��2�d&4&4&4&7�o8�q��BcBcBcBcBcBcBcBcBcBcBcBcBcBcBcBc@�@�@�y����i��8HHHHHHHN��q��\Z\a\as�s�s�s�s��9y�9y�9y�a���o��}��0�q���7�a���o��}��0�q���7�9y�9y�9y�9y�9y�9y��U��5:3�Fx���<tg���ў�oa����oa����oa�j���:3�Fx���7���{�7���z^���9{�/|��h�}�:<�]�/;TV���c��Uj���{����U�V��ԽԽ�+WV����{�WY��]h�=g���Q��3�Fy��]c���k��Y��]f��u��5�;��f��u��E�=g��h�~�3�u���Q�:���uqEqUqU�]�]�]qU����o��	��M�c�9�c�9���i��Z.�P5^e�2������6�����_��-�h�'D�tN3����8��Ф��}�[�3#tN7D�tN������}������8���8����������jK��U����'�vO��
�c�ꍸFsFsFsFhX@�PL۲�J81�l�g"�H��($�	&��}I���Ro��|
O�yK<��*�����������ǚǚǚǚ������������������ap��W�W�W�I�g'��UT�'�I�R/)��E�g������
y7�Dߑ|�
r�)ʠ�*���
r�)��O>
y�L�&�K^%�ݤ���*K�e�{d�{d�{d�y+�䯿���J����u�*�{���^�qW�~���|����l��l��l��%�^K
����������������2|<2|<2y~>�����w���XQ䯿n��݄��'r�\�W+#vůbұkص�[�-����r�\�T�(��Fϲ2}��Ռ�������������������������*�J�YX�F#���`B0!o)7���M�&�yI�Rx�'�I�U�V=V=T�
K��[�z�7��z�2�p��F\)9�I��Nw�s�������}';�3#3#tN7D�tN������|g�Ϲ�s>�}����2D�ND�ND�ND�O�de�޳����	��2�7�o8�q�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�m m<�y���4���Ӂ����������������qiqiqi�]�]�]�]�]�]�^|���^|���^|��q���7�a���o��}��0�q���7�a���o��}��0ߢ�EV��Z*�Uh��U�^|���^z*�Uh��E���<tg���ў:3�Fx���ի�WV��]Z��uj��WV��]c�<tg���ѝ��WV��]Z��uj�����~��}���o熏<4sU��ի�tgj��ի�WV����{�{�{�{�{�WV��ў:3�{��Y��Q��3�Fz(ϭ[�տ�[�(���(ϝ�;��^�{E��^�{E��^�u�������7`e��VwWW]jϭY��uqFwW]jϭY��\U\Uu�u�@�y�?6���������}��i������;�]���:�Z0��K�Z�&4&4&4&4&7�O�����8,�,��
Nk��u��2�2�B�B�BÚÚÚYvYvYvM挛�7�2o4d�h� n� n� nɼёBQ�BQ��V��Yg��o����*��������L��gg<۲�J95eT�pcnʩ(��ݳ����ʒ���_p���%�RΩ=¿B�B�B�B�B�2�2��7�B7B7B7B7B7B7B7B32327B7B7B������'������g&�;?+?,���97T����dBO"y�Ȅ�D$�!'�	<����(F�#?�?�_�	�݉nFOr1�_%}�v۰���r�nX7,���r��`�vX;,Vx�h�XѹXU�XU�XUۯ�ۯ�ݍ�r���%�+<V4nVnVy,*�XQ᯿~������'�b�rX7�'�^߯rX9,���vů`ݱnطl[�.+��bܰn�O^�z���]ό��w>
y�Sς�|�য়<�)��O���U�B2>�>�>���������������_�/���E�"��@��*�������c�p��R\).��h�h�h�������������
NjNjNk���D�D�D�D�D�D�D�D�D�D�D�D�D�D�D�AhF\) o���'�C�d��cBcBcBcy����4&4&4&4&4&4&4&4&4&4&4&4&4&4&4&4&7�o8�q���?���4�4_iiiiiiii�2����<.x\�-.-.0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�Uh��U��EV��Z*�0�˹˹˴Uh��U���<tg���ў:3�Fx���ի�WV��]Z��uj��ի�WX���<�o�V�WV��]Z��uj��ի�4Xh��a��u�^|���j�:3�uj�V:3�U����c�<uX��V,4Xh�Uc��U�^y��j����\���^|���^~p݁��^�{�՟Z��V}j�E��^�{E��^�{��:.wWWW]jϬ�^���+���+���g/;�wWgqEqE֬�՟YwYwYwYt�hL(KHKHKO�_��@˺�@ˠj��@�y�?6����?���i����&%�d��o��8љ���
L�M
L�Mkk����5�5�¾�u�U����77�2�B�BǚǚǚY��g���M�ro������F_"�K!�d"Y��I�����d"Y�B$�Ro�����,�uK:��R{�~���O�'�Яа̰̰̰椸XsR\,9�.ԗ
L��k�kjK��5T�����?���<����rn���*��B2!'���	<���I�}d}d}iB4�P�/��&�Kr2{��(���g�܍nF�c����dKV1�׍kƵ�Z�(֔k^5�܌nF8�g�>(�ܩ/�R_�;�%�*K��n�XQ߯��_W�O/�_�}��׸lg�`߱rX;k��'v�φN�o׸kܖ��vŻb�qX��\V+��r��ce��T����ύ��G>2�e�X˺��uc.��]Ռ��w#�#�#�>
y�Sς��M�Q7�}d}d}d}d}d}`�`�`�`�`}���}���}��ȿ��Rx�_�_�_�ap���ꤸR\).�ѼѺ��������ԜԜԜ�7����[�:�p��F\#.�˄e�2�p��F\#.�˄e�2���v>n�@�p�����s>�}����4������p�ИИИИИИИИИИИИИИИ�q��y����NE�/��|��������\ι�s.1�-.-9�s¸����¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸¸��.�.�.�.�.�.�.�.�j}mN�
���������4��U�5[�U�5[�U�5[�U��<tg���ў:3�Fx���ի�tg���ўj��~j��<tg���ў:3�Fx��ګ;Ugj��U���\�]�i���UX�˳K�6iy��ц���֥��ٰ�ah��i�Ӝ��������
�
ͩ���w��|%��Z�%������]�]�]�]�]�]�]�]U.����]���O2�8P5P2��8_�-O��;��+��������(HHHHHHH----��s?���U.��y����i�h���h�4��sD�O5$��3��8ޫ����O	9g��Ro�d��&�vE	|����kk�UT�,�|���˄��,�I�Rh�&�I�V�	?T�"���`}�����R�FcJ���}\Ĳ�aG>}�*��U�t������d���V~X�0����������v~V~V~R(���]g&�97Y��Rn�����g'�I��O�\+���g'�I��Y�"��E�g�x��	<Iʾߟ���)ʡ�D�����z�-x+�#'�w�2}�7{#'�>���FO�2|Q��F��I}ʒ���5���Q��߰��{���`۱qX��\V-���{n�|U�⯟|����_=�	��O~�|5�����_l��l��}�5�����K(¤�b)z�����BEv&�
�_@�]��N!,��t	5��&�"D%��2'v�*�ʽr�\�ܖK%��^ۯqW�v����[�T�s�j���ױ�װ��aG^��{
:�u�(�F2#������J��*K��/׍�^6�x���o׍�^6�x���oό��w>2�|e܈�9�r#(�FQ���
�+�`���<��������&�97��<���a;�@��v3����� ga;�@�ǪǪǪ�v3�������a;�@��v3����� gIp��R\).�
K�%���v>n�@�p�����pZ'�pZ'�p�/��|&��4_	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	���7�����NE�/���o8�q��y����4�4�\ι�s.1�1�-.-.-.-.-.-.0�0�-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.- sN4��u��qiqiq��^y�ߚ���ߚ���ߚ���ߎ��ў:3�Fx���<tgj��<tg����ߚ��%��~j��~j��~j��~j�㗞9y㗞9y��i��cc�a��Ej]�5�l-�-4cs�>y��1�f�э�F7<�y��.1�1�1��u���2D�ND��}���	�	�	�	�	�	�	�	�	�	�.����O���?�y�@ˠe�2�8_�!1��s�����\Uu����7��Hhhho��>o�����$� g���XBU��/_�^O��&�|M�<f9<f:����e�����U��/_VO����Ye�l��'�2��e\�|L2�9�8s�p���Ұ��akJ�֭~=Z�y�8s�p�XZկǯ'ͯ'��,��'翁�����;���|�����Չ�k���i-�V4�=7~Ye�Y%���=��&�V�w���ζ���SuKow-�)G�R6EX߰�n}�`�ғ���I��Q)T�"oό��G"&�W��_oȂ��vU����pa/����K�>��������a/��<�`����_��r��e_o����$�PS�}�U=(���Y�SςiD߫=���i'�Iwr���K��7�R]ܱ�r������w,o䰣�_~�}^e�eT��BE/������@����
�]�H��I��ɮ�0p�0p�0-D0-D0-~`ڈ`Z�`����p*�l���2�|1�V����BMF!"�@�U��U��ڶ�Z�df�g����pe�2��
��
�{:1{:1{:1{;��w�dS�ȧ@�(eD�H������{~��'o�������|�yܤ���]װ��cwJ���%^�����{+��W�쯫�_W���e}\���R_�I~�%��7uln���ձ��aWr®�]�
��w,*�XUܰ��GJ6��m(�9�s�j���ύ��I/�I/�W>6�|m\��815pbj�AQ���g��۲o�e��e��e��e��e��e��e��e��e��e��e��l ga;�@ο���o���'�v�v3����� ga;�@Β�Ip��R\).�
K�%�'�7��|ݱ�v2���q<��|O;�y�������w�;�y݄ƄƄƄƄƄƄƄƄƄƄƄƄƄƄƄ���4���ӄ�|&��4_	�����4�������O�i����~n:::s:�u����7\n��q�ڟ[S�����������������������������������7\n��q��u���:/��8����7[S�/<�o�V��o�V��o�V��o�Fx���<tg���ў:3�Fx���<�o�V��tK��V��o�V��o�V��o�V��o�/<r��/<r󱍸эV��B�6��B��Ƈ^w��>����}y�ל��9��@�@�@�@�@�����B������`o��v7���<ݤ�v��J��e�����ȣsK"mI�ɣ1�X�ȓ��I�eU�t����r$�9x�<�������-�+�Tg&��7���O�,�فߕS�;8u�Z�(��M�Y7od��^M��"�ϯ׳�*��aq�"�ܕFnJ�7ePR�����Rk��>�x6�,1ʤ�$Ѷ��sJ��R/:�.-ZNM����?&��ޭ'|f�G�̈�̏�,�+�|��m�K���[;�y7>����#�r6��݌�vD»"b�����m�����_XߓӸe��eo�MM��S$V^�;/m����A�H<2*n����&���+|�z���o�O[߰��I�{���
��;�·
����,D����\��^,��ْ�`H1	enc䍅ny����gW>���zT�Ҥ�J��*K��h�R_�GJ6��m(�:Q�s�.���ω��w"
�D܈��bh��]׌��G^2��m��}ZJ������wi0�����a�ù'��&��,͹,��a����ܲ�m�
�)d���7䫜7?�7K�" ��7���ߘ6�03~`������k�E/�gVg��/@������pp�pe��0��{;��6��{n|�7�*Ew�M���N��[׸�`�YՆ�����بk�..���H�M*�I����킐�.2ߑ2��vD�[�6��jۑj�*�Mո�8�1|^kz�1|^r���A츦�f�jڬia�����*��*�,�Ӵ�Su��,��F; ��eo�7���e�)=���챿>6y��ƭ��[��.�RO"1��D�#�7��߫c~����=^)6�<|��,*�XUݱ��Iw^6�x���.��]�����ǻ'ͫc�"2����>m*I}*I}*I}*I}*I}*I|��9�eQ���yTd��2_2�e��X���p��᳉�g��'�N8�6q8e��e��e��e��e��e��e��e��k��_���7�������o��}�� ga;�@��v3�����z�7��z�2�p��Ah����'��Z'��O�i��?��	�	�	�	�	�	�	�	��4������sO�i��?���4�������O�i��?����7�o8�q��y�����?�_	��'[��/��~y�4�sN4�sN4�sN�8��8Ӂ�8Ӂ�8Ӂ�8����7\n��q��uƸ�����������������8(y<o\d�&}�n�
����З����<4sU���֮�]Z��uj��ի�WV��]Z��uj��ի�WXoa����oa�����R�R�R�Un��Q��W��h�������o�G���������4��ϗ�/>^|��y�B@�c0��a��ږRc�X�Xh���'��������������*�ݕAndD�dD�qK6�i;0~��BndD��XD6�P��U�M
�I�W)4*�&�\�Ы��r�B�Rm���4���4�'&��V��$j55�G+c����[���{y���1=�[�1<Y��(L��zR/=�?weP]�?�T�l�e�k�Y��ɣh�#.�#hȬe����hɣe�,1�ɹ��@����ȉȖs�I�`�泱�gcj���}�T�f���D�6�U��|�֬�7e�=�<ۖy�dX�$ֻ$ַdX�,�nY�ȱ��cw>�}]*���y}Y<����&�TM�TM�0S����`����aGV��[
:�ul(���կ��^��`R2+ڲk��*9�
Ge�]yyY5�)e��y���^��J�R���%*�J�R���%�������`B,������য়<�)�Dߥ~�e�X˺��r>�>�>�য়=(���o҉�E��Ҥ�^���[��w+�ʾ��Z����r˻r˷)=�U�⯟|����_>*��Wϊ�|U��ϒO=�e����$��I���_�"V4��eWb����ȫmϗ��U�ʨ�pe��1yU��Bά^Uj?��?��?*Ë��%o�H[�2�#�3+�e��(\��[�R��_��Ri�#r��/&�E��]_E�WY�exi4Ы4*�Jጶ���c�ʭCpe�btaR+����5�K݊!"�N���a�I��#��XƔK"	*�������dF4�'���`}J�Y�TK	����������D���YR�F����E�'ǟF�&�Y�$_����E�"��H��_��)g���Y�,�yW������o��}�U�U�U�U�U�U�U�U�� ga;�@��v3����� ga;�@��v3����� ga;�@��v3���oY���oY�\#.�-��8�w��D�O�i��?���4�1�1�1�1�1�1�1�1������sO�i��?���4�������O�i��?���4�������O�i��?���4��sƸ���2���;N��q��u�������>��q��u����7\n��q��u����7\k�K�K�K�K�K�K�K�NxP9���X�Lt�sF�c�����W�j�q���GD��tgj��y�]Z��uj��ի�WV��]Z��uj��ի�WV����{�7���{�7������W�诰�qp����~`g����������������������HD$"��AB �17lbn�FQ���_VOI/,��,��a�����]���'��'��'��,��*��Ra��}'��$�>�a��I��U����#0ɣmK#0��U����x,>ь�F���hH�3ґy�ұ������gY���&��I��+�����y� Q�Q�+�<L呗��gc����XAN7��c�_}|mYe�5��~;��}���7�7�7��c�RU�Fѓ�ξ	,�H�/���*�����2�8�Ƞ�(%�L�#/���O�,�K!�D��M�"�H��1�pcn�������w6�m�۲�D�,�K!�D�,��}iK/�X,�X�U�"��^�X+��dM�F,�X�K%���`A0 �L$��E�"��yI���)d
M�B%P�T##�#�#�>
y�S�������B%P�T##�#�E��հ��'�쯫�cw>5����D�c]�7���v�{��ݯ��|�k�_=�����v�|U�*�ܲ��e�2k�2k�2+�l���݅Y�?�V��8T�
�(�pn�p*�,���Xiں)ڼ�8$R�q|��Vj�nF���k�Ov��ַ�׶OvA��Mׁ��h��!+z�i��:��r��Y���XYwi9,*��o���XU��D,�D,�B�X�R,�k]��<2y~<�7�l��cK�K�r1�,�/*��^ۯqWϊ�{�w+��W�쯫�����`�%Q)TJUȌj�ߥI<����g��dF2"oȉ�U9T�>���>���>����U�Vkj��}�ǚǚǚǚǚǚ7�7�7�7�7�7�7�7�''''''''7B7B7B7B7B7B7B7B7��z�7��z�7��z�7��z�2�p��F\#.�˄e�7��z�2�p��D�Ah����'��Z'��O�i��?��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	���7�o8�q��y���4�������O�i��?������g\θ�q�-9�u�����ڟ[S�j}mO����>�����ڟ[S�j}mO���a\a\a\a\a\a\a\af�ͅ�6l,�Y��af�ͅ��E�l+UXh���U���]Z��{�7��uj��ի�WV��]Z��uj��ի�WV��]Z��{�7���{�7�ޗ�����������iת67�,x�����@��`P0(
�HD$"��AB ��_`_`P^P^Q?�?�?�0�����$�a'c	;I�}����W�)<M���k���x�1�(+�d
���0�i?�p�q.��27�员la.���E�������O���BhR�2�p�������'��"����������F�FB#!�g�v0�i?�|�2������������I���Dݑ}����Љg���M�}����"n�D�����w&�M���7dЉ4"E�r/��}��	"�92���#/��`F_���`F��I4J�1�bϯ��&��&�בQ��`R,�(Ě	,�K>����FDl�#g�<�˹�r#.�F]����Y�,�/���M�"�H��P)������#������	9T�_o�AO�"2�%\�K�PS��Y�0>�Q)TKJ%�I>��,o챿v��e���7�X��ce�����vŻb�X�V��n��^ۓ����c�N�!Vs��_�^�R7bZ_[��J���g����WхJ����ߑs��%X�nG�Ƭe�;����mX˽��eP��)��3vF����ߑBp��Ռǥ/�&��"�Սå/�/�G>&�D܈+���ʾ�*�ݱ��Y��J��I�ܩ/܌qR7#]��x�|K>%�����װ���'�yg��V��OՑ��`}H���Ro)7���������E�"��H��_ԙ����1zM+v
����Ωd
�����������c�c�c�c�c�c�c�c����������������������������������q�˄e�'�'�D��D�'��Z'��O�i��?��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	���7�o8�q��y��	��M�h�E�/��|&��4_���N�~���G�Z�zՄ����ۋK�K�+�+�+�+�+�+�+�+�+�+�+�+�+�.r�r�r�r�r�r�r�r��Y��af�ͅ�6l+����<�V���a��E��^iy���z�ի�WV��]Z��uj��ի�WV��]Z��uj��ի�WV����{�7���{�7������h̗�͍��VlhO����������������������?�g������3��|�����O���3�����}'��?�I��'�4�h�}�I��'�4�h�}���T�6֮�M��)e�^ǳ"&��3��D�ǜ��E��7~�#<��p���C��'4o�2h�u�`j�u�'��,�����޳���7��zΒ�ިިޫ7�BN7��a�c��FuF@�|� Q�(�d

���Wޫ�i?�|d
2���'�O4M�3�2c���NO	9g����������NY��������������+*N�N�N��
���ʿ�O��$��?Ԟ'���I��.xFc>��}\���7piU�s���X���YĤ�I?��e���F_�~M���7p"n�?����)<
O��������	?T��,�K:��Rh��M�yH��_�/+8E����+�U�+�K���}���FM�&��yH���XX0K8E�"�g��Y�0a0��D��#�#�>	���ܱqX;e��`ՠda���r�k�+}�x���av?��/��r¬K���r�Y�j����(��/�ok���N}�V����/�9�=�Vx1��d~����ϖo���eRȆ�_rU�ȶܳ�ܚ��.�ŋ�qb�RCrB�nHQ�
!�r�}�����X�j���s줫�p��⯗ܰ��IwV2r�)��Y�$7nG�{;���������U~��{:�2�T�t�*�����a쯵�I/�I/�I/�I/��"7Dn��6n�dFV�r-���/��J2�J2�Rx�'�I�V3����� ga��H� o�����H� o���������}';�9�I��Nw�s�������}';�9�I��Nw�s�3�g�Ϲ�s>�}����3�g�Ϲ�s>�}���p��F\"y�y��>�}̉�|O;�ND�������N�7�o8�q��y����i��?���4�������O�Z�zՂ����&�\?n%��K�s�s��9y�9y�9y�9y�9y�9y�9y��U��EV��Z*�Uc��Uj��U��UV��Uh�w6�Ua��Ej�6�Z���֮�ў:3�V��o�/v�ի�WV��]Z��uj��ի�WV��]Z��uj��7���{�7���z^���9{�/|��7{+�7d��������o�p�	G�%��~�Q�	G�%��~�Q�����W���_�����8.���8.���8γ��8γ��3�d47[N��m<�@�@�BsFy�c�^��$%_������.�~�_�C���$&�>s9˴Us�@����qu�n�_��Ru�"��U���g�����!1��)<��!'c�����|OTOTM�&���������֌gY������h˄O4O4e�6c�c���걸�'4n�n�'5���n'cq;���N����7B7B7B�����h�!(ɾՓ}�"���DѰ������������������"Ưd�6�=yf9U%Y���2�8����E�A$PI7Գ�Y�,�yK<��R�)g���ǚǚǚ�B�B�272ǚ7���Ip��X�W�X�RhFhX�F�X�R\,.
�������Mό���@׌�����?�!�?Y7�D߁��``B0!�T"U҉iD�#'�>����Ov6��I�X.Ry�Ȩ�21�t�vʱ�K.�F5��Xn���~�8��rk��7~�J��*2܎�8�σ �#���dR�!��\q��LRG�3�b�A�ҳ���w�)��W=/K�H���yY���us���#��)�r�?���W����K+1^�VH��Vb�,���,��zYY#�M��O��i�}�LyV�,.8p?ܥ����7+�n��פßG"2�De��N�6%��v�P<2���8��R�*2���?n��_���&�DM\�ڶp�8F�Ⱦ�E	}�۶n���&�VM����Y��
^E/g��'����ap��R\).�
K�e�2�p��F\#.�˄fdfdfdfdfdfdfdfe�����7ln.��]���cqv6��g�Ϲ�s>�}����3�g�Ϲ�s>�}����22�p���Ђ����2'��<��8-���O�i��8LhLhLhLhLhLhLhLo���?���i�����HHHHHHHHO8�q��y����7�n��9��E��������`q����Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��X��a��E��,4Xh��a������Ej�6�Z����ў:3�V��o�/wD���m]Z��uj��ի�WV��]Z��uj��ի�WV����{�7���{�7��r����~L�L����c����Ƈ��|����=n��w�[�z������������s<�y�������O���j��щ����ۋ��_	�p���^��9�m:�\ah��E�4�������O�i��?��Ϋ�i�@���c���'����ӱ�/���g�������tg;�s_cVO	jO	j��$�e��e�zΒv>o���e�'�&���s �N��9���9�'��-��p�ИИ�q��"tN2�p��RsF�FfD�D�dg�o��Y�Y�:'cV��'Z1�cn.�s�3��:'	.��i���I�Ip���'�vO����?��xI��ݓ�NǚY��w&�ʓ�7B��E�r/��}����_g"�9�ȡ/��򰁝�� ga;�@Γ�7B7B7B323232327B'�7B2�I��v7��8��-�Ȟh�˅'5'4��Yd%?�l����ëa�o��f�n��yT+�~ݕD�Ҍ��I�"2�De����s�h���ω��wr���<U����qW�ܤ��R|<R˻��ݯ�������_������D�
z��y0 d�<�Z�[)��#�l�$�G+eo����t�t,����`�_�������d/��~�ms��1\��[��gK�B�-%o/P:?��!f)���Sǅ���I|�K���k��mw�����o+�7���o+�7�G񷐲VJ��s��֣Z����Γ"'�|n���ZQ�t�p�RK��Zϱåc�J�54��Y�,�I�R(�^R���?n��"�u��&�9��'�K<��Ro�e��e��e��eT���j���e��l|ݤ��%�Ip��R\).�˄e�2����w��'��<��|fdfdfdfdfdfdfdfe';�9�I��Nw�s�������|N��h���h���h���h��Ϲ�s>�}����3�dO4O4O4O4��&4&4O;�y��pZ'�4������p�ИИИИИИИ��?���i�����O��6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�*�Us�\a\as�h��U��EV��Z(�E�=g��EV��Z*�Uh��U��5j,�Y��Qf��E���UZ��Uj��U��UF��Z��Uj�����UX���<tg���ў:3�Fv��]Z��uj��ի�WV��]Z��uj��ի�WXoa����oa������^���9{�V�5��v��������j��ǅ�<,xX��h�э��F6�M�W��Q����|�5��������5�9��㿭��as�s�s�a�٨�q�	ά':�mO5�7`e��Vw]j����Q��w�����f�����5޲�sh./}�F��ۉ2�^e�&��}�?�����W�h�h޳���7��y�� ��n��BcBc�?��	��M�\Q��|���Bc}����q:'��˄e�7B'��tf��8��Z���H,s��|f�����h���Nk����HL(�����}���:�_vO挳�[�������z���q�V=V=U��h+���15l�ճ�w"7d��Dn�IyTm\��nȡ/�����|%d%d%d%%%%��7�<�,�}�[�:�cqv6��m�؝��8���|g;�n.��]���cqv6��'Z4�h�u�cV���[�� n� n���I��cq:��o4e�7k��y�y����o��'�vO����?��o�d��ɿݓ����~n�����%�?n����e}�۲/�d
E��9Tm\��6<ݒ~������]����b�X��fFF�Uٯ��Ź�ɷ�ɷ�r����g����nB��!]��=��wf������o7�K�MI*�X����`I��n>�y���	�'�$g�Hȟ񑐑��b`���y�'��ϯ�����ϕv�ʸs�P�,���>���N�אb�6�(E��(�n���
����$�wm��M���S�w��n�B������%[w�m�@␢�CrJ���U��J����rIT�ܭo�M�b)��wn��ܭ·7l�+��\]��]c�폛���c���7������7i o���7�޴czэ�F7�޴ln.��]���cqv�������7c3#3#3 �#3 �#3 � �ND�ND�ND�ND��}����3�g�Ϲ�s �N�'����LhLh�w��D�O�i��?���4��yƄ��	���7�HO��6�� m?�@�@�\Z@�\Z@�\Z@�\Zu����\.x]p��h��U�]q�q��]��EVj,�Y��Qf��u��5�j,�Y��Qf��E��5j,�Y��Qf��E�����*4Th��Q��EF�^]��Z�ի�Z�^]V�^��Yګ<tg���Խ��oZ��Ej���4V���Z��Ej���4V���a�/u������XoK�K�9{�/|���R�xV��j�K�c�^tq�a��Uj]��5��t��5Xh��a��U��V,5Xh��a��U��iy旞�7��~�7旞:�TX��c��U��V:�tg���_~k��}���]f��Eέ���q������;�.r�r��Fz(�E�=g�����^�8n��?2��KS��}��zH�z� Q�gI�����W��r�r�/9�q������C����9�8��!1�1�1�1��}��i���L7a0݄�8LhLhLhLh���8��̂�?��6�6����}'5%�3�3�3�2�c��l��h�u�e�
�����c���7��X�Y��g�����&�d#6�Td��%¾
�'���g'�`B$�Z�2��2���d�j�����	�a�&������d�8`���j�UFfFfRsX�I}'��(�v�:���ԝh���/qF'��ˊ68e���Q��l`eR�L�7�+8�+8�+8�+8�yN��'^E�"��v`B�0!]���Wf+�ف
����vV?4�ߚU���oD~UߕE��()TV�
�Sh��ݿ˖��F�Mgg�"�����Օk�ikܵu��wy5�73�a����������-��s??��^����*��Յp��8���ݶ?����r�����̖�;%er�lF����l��/��c������3Q����QH�����!�˜��K�6�lWy��}��s����������r���g2_�=�
F�!Ҿ"��Y\~�����v�>�R�!��4R)���u:�>�o��(px������=�>�ƹǷ�M��S��a�\z���krغnJ���q�,_�?��֌l��7���I|l�7���p��D�"n7��M�&�����������������pZ'��-�h�E�Z/��|�������sO�i��?���2�d&7��Lo9�s<�����C�����?��8����5Ť�Ť�����WZ-.0�Z\ah����i�]���69vl.r��Y��^y��^y��^y��^y��^y�玫V:�TV��ў:3�Fx���<tg���]Z��uj��ի�WV����������U����Vv���Yګ;Ugj���U��EV�Z,4Uh��U��EV�Z,4Uh���K�Q����u/uF�^�Խ��{�7R�R�R��^���9{熋��a���Uc���Wz��/<4Xh�Uf�~l7ڪ���UV��UZ��Uj��U��UV��UZ��Uj��U��/~9{�a����n㗾�YᢵVv���Yګ;Ugj��U����v����}��ߚ��]f��uέ���q�������0�˹˱ў:7qѻ���ў:3�Fz(�E�a���p��V}j�����������&���:O��@��P/��m.0�q��y�|i�����C����9�8�8ИИИИ�m>�}���?8n��v�KS�ƄƄƄƉ�8���8,�,϶�6�6��'�q���7��M�'�6�γ�����-������BB2�p�ƌ̓��Y�*��'���}`�Q�}�Ǫ'����x˸�d�V	d�5�_:oLC?���'�ЁD��v���7��e��j��m���p�fXu���oY�\>�BfF\,4__���E���Eo}r/�r�r��.Vw/��l69�F�S���6�V����򤭏*J�򤭏*J�򤭏*J��$�n������\^�J��2����(l��Ce%J)+��m��6)Sa��n�)S��:!(V!R�b�ݬD7��BB�V$*ub����!\;�������7�/�P)ШU6
�b	@�V$+om:�@��쏑��%l��@!�>�����uG���!��>����C�<���v
�7���)��~?��U�-n/m�,����Ch��T+~!۷
����������������������չvirk�qFD�ɤ�l��,�	<lll��Y����,�`�$�5�k;
�%|���Ec,���RX�),dV2+:�	=~��O_ş����������۹����m�y5�zэ��6���`o���6���n7��M�&�p��F\#3#3#3#3 � � � �"y�y������������NE�Z/��|��_��-�h��i��?���4������sO�g��9�s<�y���3�����?�����B4�sO�7\n�����WWWWo��}��0ߢ�E��M�-4Zh��i�6l,�Y��af�ͅ�^y��^y��^y��^y��^y��^x��c��Ej��<tg���ў:3�Fx���ի�WV��]Z��uj�^�^�^�^�^�^�^�^��Yګ;Ugj��U����Vv�έZ*�Uh��U��EV��Z*�Uh��U��EV����7Tn��Q��uF���7Tn��Q��uF�^���9{�/|�Uf�<ttZ������޺%���+UY�ߛ�����a��E��,4Xh��a��E��,4Xh��ߎ^��n��w6���Vxh�U����Vv���Yګ;Ugj��]����]����]��ի�TX�K�F��<sэ����<tg���ў:�Z*�U\au�>���]�]���3]����p\�7��<݂�B\ �_��q�q��Bh�E��NBBBC�g\�HO8�q��yƄƄƄ�8KS�j~mOͩ����22������o��q���2BBBC�7���O;�_�pZ'�C�7�ho�Z'�3�4�'4������h�j��4��czΒvq�wptr`�ȌK.P�Y-��E�WY���ZςI�Q��o�I�݄AK�!(�\)4 h��p�@�O��|%�3���C�46;?8��0��K�\c��E��������8-��Z����n1�玎,4Xh��a��Ej���R���a0�J������f�5Y��Vj3Q����L�2�v�uLf�A���⊎�s��F�k�~�U=�iR>=C��e�u*H�S�j�kQ�l$:fN[�֪y]6����d��uK�L��v�վuf���nݻv��h�V��f�������9ݚ�D�U0�L&	T�Q(�J%�T�a��l<��熎j�㺌���q�g�q�g�q�g�q�˄e�2�p��F\#.�'�q�'�q:'�q:'�q:'�pZ'�pZ'�pZ'�pZ/��|��_��-�h�E�sO�i��?���4������~s<�y���3�g��9��?�����C����9��}q��uƸ������¸¸¸¸�}��0�q���-4Zh��i��E��L�Y��af�ͅ�6l,���/<���/<���/<���/<���/<���U��U�+TX���<tg���ў:3�Fv��]Z��uj��ի�WR�R�R�R�R�R�R�R�V���Yګ;Ugj��U����Vuh��U��EV��Z*�Uh��U��EV��Z*�Tn��Q��uF���7Tn��Q��uF���7R��^���9{�^z-]��V�5]���~�Wn3U�/<4Xh�Uf�~l7ڪ���E��,4Xh��a��E��,4Xh��a��/~9{�a����n㗾�YᢵVv���Yګ;Ugj��U����v�Wo�v�WV��]Z��E��4��Zh�э�5�9v:�tg���ў:�uZ*�Uh����j}mO����ͩ�h�7�X�w�h�M�6�O7b|��T%�·[Ho8К/��p6�::::s:�@�@�y����4&4&4%���?6����ڟ�o8�s!1�3 ���\�t �>�}��i����o��s>�BfBfAh��Ϲ��4��}������dL�<���qv3����o�i:�n0)g���ձ�}�Y7ڻ�|t�H�o$Nܲ��'�M�#ew$��ݻ����exi!X:0����)TM�o,��5�	d^�ԛ�Y�*��a�c����	�cvO���?[Q8���>wR�U*�.��v�;��9ښ�Fj3Q���f�5R��J���WV��j����j���߆��n�v��h��U��E���\r���玮iz�j՗�F�۷nݫ}Wh�v��h�՟�7��F'�,�v;l�~�++:<VVtp~7C<��P���և!Ԣ��uv���nv�n= �9.�?F<2��㽚��UZ�7�^�r��Z͢_:�jޗ����.�U/EV�[��熋����wT���Y��(�՜��p��j���tK��/wD���y��v��w����U��f�6�y�p��F\#.�˄e�2�p��F\#.�˄e�7D�tN7D�tN'D�tN'D�tN'D�tND�ND�ND�NE�Z/��|��_��-�h��i��?���4������sO�g��9�s<�y���3�����?�����B4�sO�7\n�����WWWWo��}��0ߢ�E��M�-4Zh��i�6l,�Y��af�ͅ�^y��^y��^y��^y��^y��^x��c��Ej��<tg���ў:3�Fx���ի�WV��]Z��uj�^�^�^�^�^�^�^�^��Yګ;Ugj��U����Vv�έZ*�Uh��U��EV��Z*�Uh��U��EV����7Tn��Q��uF���7Tn��Q��uF�^���9{�/|���E��tK��/��o͆��㗞,4V��a�6�UK�a��E��,4Xh��a��E��,4Xh��f�~j�藻�^�{��ߎ��]c�<tg���ў:3�Fx��ں�uj��ի�TV��Qc�c�f��i��6<,r�UV��UZ��U����EU�\n����u������s��Ns���3�ؘ�� q��\au�����]�w'q�w'��5ťŧ[S�j~mOͩ��?6����ڟ�7zڟ�S���g��9�\�\�\�t>�Bc}��i	jp��	�	�	�	�	�	��4���w��?��t>�A\:�Fy��~p�.*��N4�
^6�I�'�H�n���7�3��j�H�gb��؅��T�!k��ӥ���BC�qG��^�O����h��]��o���{r˽�l�[r˼�v~/~ǒEj?�"�XsY�_c��XANO/'�/I��$�������V�tg���_~k��Y��]a��Ej��Vj+UY��Qf��E��5k��Y��]f��uFk�j3Q�����^�6��Vj�R�D�a1���U�߸p�Q��&B��ht=��k���X1#�>s��;g��]��q�*��e-��DV����r�n;C��-���w�q��c��h-��ujkE�	��Ɖ挸X�R\).<�m:�}������ q��ЄƄƄƄ�����4&7�Ӂ�>��q��u���7�(xM�ZBh�6|�O��y����w�s�3����|g;�9����w�s�3����|g;�tN7D�tN7D�tN'D�tN'D�tN'D�ND�ND�ND�ND�ND�ND�ND��}����3�g�Ϲ�s<�y���3�g��9�s?�����C����� sN4��u��qiqiqiq�q�q�q�q���7�a���-4Zh��i��E��M���af�ͅ�6l,�Y��^y��^y��^y��^y��^y�玫V:�TV��ў:3�Fx���<tg���]Z��uj��ի�WV����������U����Vv���Yګ;Ugj���U��EV��Z*�Uh��U��EV��Z*�Uh��Q��uF���7Tn��Q��uF���7Tn��r���V�Wz��_�:8��j��V9y��Ej�6�a��T��,4Xh��a��E��,4Xh��a��E��j��~�{�%�藻�������:3�Fx���<tg���ѝ��WV��]Z��Ej���,r��Y��af��.�Uj��U��UX��c�c�h������<.��t_	�����3��Y�y�|Y��u��i��C�i��s���;���;������ӭ���?6����ڟ�o6����ڻ���6�����y���2������Lo��m!0݄�8KS�ƄƄ̄Ƅ���sO�;�_�p\ї���V0�`� e�h��Aa`AQ��I��cnʩ(��}�AZY�(u���6&�*�K�_���IR��C�\����5f��CiYn-Ol��փ����m�ʛ&����$)T1!�a��\����gxxe�t���_���K<� V0)TN94��K�+W�ޫ5Y��c��E��EVl-�1�m q�m q�m m m m:˺�u�u�u�u�u�>r��F�9���v5߼�����5_�1��_֭��������,���&�>�v��,��H�w$R�?�ȿ_)#K{^7#�?9�%l>��VkQ�}*$S�2D�C�V��쥳)���}��S/]����ď�l�Y+<��LO��5{%��l!3�!5�c8���rnK97��r��iTe�ZKZ��l1���ݰ��_��
vv6���}(�y<�l�D�E�e[8ʲ(�2h+�(K�P�ɿ�O	9?ڵ�Uk���}�a	V���lѯ�/_�^��γ��v��gY��F�]���qv6��m��ۋ��cn.�s�3����|g;�9����w�s�������|g;�9����w��N��h���h���h���h���h���h���h�������3�g�Ϲ�s>�y���3�g��9�s<�����C�����?�@�i�����������
�
�
�
��o��}��Zh��i��E��M�-3af�ͅ�6l,�Y��K�4��K�4��K�4��K�4��K�4��K�V:�uV��Qc�<tg���ў:3�Fx��ں�uj��ի�WV��]K�K�K�K�K�K�K�K�Z�;Ugj��U����Vv���Yբ�EV��Z*�Uh��U��EV��Z*�Uh��Q��uF���7Tn��Q��uF���7Tn��K�9{�/|���֝y��Ώ<�ڗK�K�c��U��Ի5�kKR�{�4Xh��a��E��,4Xh��a��E��,���/=oц�o�/<uV���c��U��V:�uX��a��E��,4Xh��Z��U�^x��j��V+UV��V:�uX��c��Uq����ڟ9w9w\o:/��~q�q��Au�g���g��	���&��q�~�u���;���;��������7�o8�q��y���ͩ��wͩ��?8�q�1�1��ND�tN23�7�O��mQ���+W�fAfAhAhAfAc�9��'5���;�(�Iy<
73>2^����7k�k�Q�a��ѷg��6��3V	!k��J}�:';�GX�������&�\d�=m�ݨ���j��X�%,D^'���v�zǣ���n{���f��÷�-Gi�T��^�����ӰsH�^M�/�/*�쌞|�+�J�%����@�7�H�5���y�����/�^7��$&ϵ`�Ռ�VM��2��N8ʶq8l�pɢpɢp�Rh��́I��F&�
M����Y��Y�"qʢq�F�ՍͫIkJ&ֽ%���I7��/�Tl+"��>ǒUc��a
Ұ����jv���J/Żɥٽ�z#�=����C?��T�u2��bk�:�'���)��tvn�!�L�OQݐ��t����rE����T�^Yc&�ͥc���7N���7�EI�&�۰�쌁���^df�L;�2���u�oՌ����J�/ү��_W"6x1,���XݕF0bX1,�	����A$PI�ɾ�����+(KK���<�:�`T�Q�Ԑ7�@�I}$��7�@�I}$�˄e�2�p��F\#.���}';�9����w�s�3��:'�pZ'�pZ'�pZ'�pZ'�pZ'�pZ'�pZ'�s>�}����3�g�Ϲ�s<�y���3�g��9��?�����C����9��}q��uƸ������¸¸¸¸�}��0�q���-4Zh��i��E��L�Y��af�ͅ�6l,���/<���/<���/<���/<���/<���U��U�+TX���<tg���ў:3�Fv��]Z��uj��ի�WR�R�R�R�R�R�R�R�V���Yګ;Ugj��U����Vuh��U��EV��Z*�Uh��U��EV��Z*�Tn��Q��uF���7Tn��Q��uF���7R��^���9{�/E���E޼���;R�Un��a��Uj]��5��t�,4Xh��a��E��,4Xh��a��E��iy旞�7��~�7旞:�TX��c��U��V:�uXh��a��E��,4Xh��Z��/<r�ڪ�E���Yګ<uX��c��U��EU�[S�j|����q���i��@�Ђ�8����2���I���J60�c.��:9����e�47��9�s<�Bfȳ��	��22B'�'�'�B33�dN7�h+W�Z�� � �#4#3#3#tN7D�9����)?��g��������"�r��������[����[���_~���~����]�Y�e
OlC5S�\b{q\Onq$E�Y���~���*A�*y[f�Wa��벇����o�-���}o8�V3��o9�Ӻ:���}1;NH�⟦�$�7���e�����g����Q�*O��K���pk����Xs��сa���Ԛ�Ԋ�_6�|m��9�s�hʩ(ʣjʣj���X�ϱ�*��*��*��*��*���I�>�6��>�ە�.U����7���e�;d��1|��|��|���O�?�ro��(NI'���8��
N
�+;>�ͺ��H�ÿU(<��Ԥu>[���(u8��Z�VkQ�պ]��봨=k'C��%����n��=���V�S��+7,6N��n�>4l���
��c���H�xd�W+��λ�k��;�����*K�#0L�K1�Ȍ`�0>�Q)TJUȌgƳ�ZT�Ҥ��1���`A,��P�d"O��&�۫��^VOj��'��A_a:H� o�����H� o���2�p��F\#.�˄e�����}';�9����w�s�'D�tND�ND�ND�ND�ND�ND�ND�O�g�Ϲ�s>�}����3�g��9�s<�y���3�����?�����B4�sO�7\n�����WWWWo��}��0ߢ�E��M�-4Zh��i�6l,�Y��af�ͅ�^y��^y��^y��^y��^y��^x��c��Ej��<tg���ў:3�Fx���ի�WV��]Z��uj�^�^�^�^�^�^�^�^��Yګ;Ugj��U����Vv�έZ*�Uh��U��EV��Z*�Uh��U��EV����7Tn��Q��uF���7Tn��Q��uF�^���9{�/|���f�ю|�_���Z�U����.�i��Ժ^��Խ�TY���0ߚ^v���c��U��V:�uX��Z��.ͅ�6l,r�UXh�UZ��.ͅ��E�;WsU�5[�U�5[�U�5[�U�5[��u���������ў�{��ߎ��]f��U�^wo�E���`p�*�ڜ&k��O�7�ˋ��n�BU��F���V���간�&:L5�o�Ɖ����dL�j�����|gY��}���	����'�
�I:�J6?�W+�'�mgF6�_��*�i��iI�&�VO	8,țJ��k�&��6|m��m�V;ogZo7��7V�B܁��ѠH�V��v�[[���#a�i65�5���ۤ�����=��\���^�^�\���~Vd�d~�o���'����tv�����l)$P*>/�ۡ�v?���}>�#��1Z�jjB�씷e���]�=+-+)��v��n���\4�6�~B�׍�J��O4N��5;�rM�32Y��I/a�����,��_G�U���偎Uհ��I~E�ݻ;�7Ԋ	å	�"ѹg�rY�
���^&����E��6����]ʒA݉��BV�#a����}}(�n�oe�=��ە��Nk/&��$Ndg++���p7����e=��q]�RH�e�4=D�l�bk��m+��e�T���ݳ��ڙ+a���>Z̞'gY��k;ܮJ�&��yv���J���`�l3iDڈJ�)۲(VE'�3rM�rEq*���������"���C^�"��av�"�ßqr�ǫ_w"�a�gҰ�V��}��)��x��iX_g�B0c�ԋ��Y�A8t�8�P2(��K+}~8�jK��U����a;��X�X�X�X�X�X�X�X�RsRsRsRsF\#.�˄oY���M����&d&d��h���h���h���h��Ϲ�s>�}����3�d'9�s�'9�s�'9�s�'9�s����?�����C��i��i��\n����WWWWo��}��0ߢ�E��M�-4Zh��i�6l,�Y��af�ͅ�^y��^y��^y��^y�玫V:�uX��c��U���ў:3�Fx���<tg���ў:3�Fx���<tg��,4Xh��a��E��,4Xh��a��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EF���7Tn��Q��u/|��r�Xj��h�=���u[�5V�٭3Zc��U/E��Viy�w����玫ժ+TX��c��U����l-�-3Zc�cµUj]�]�6�m���V:�uX�ў:�tg�����Fy�ߎ��7�^kWo�V��sK�E��U�����0�]y�8L�z�\Uy����8�s ��n�gc	vOvYvMvO9?�|"�&zU�t��Ⱦ�6�I?�К���F7��:�`T�Q�Q�(�h�h˄e�7��a�gw>Y/�'�"�K �(Ŝk��"���h��}��`F,�ݤб�F�Ҥ�,��dF]դ��v���BEܓ���X�� �Z��h�t��eS�m��p���K�Z�m;�	��X�rV:nL1
�/J�(I�K:��MK���=_�����qI}F�s���ۖq#B�f'�8�B�dv/s�`TrT��S���;|	#���!PbH�x5�o�$E�
d��V$�wMs��mv�=,���m؉Y���+r��$,�#�c[܂���ȌY�p���u�uc.�y`B,���/���r�Ƿ"������"��_<���jUձ�Mհ���F7,�g�Qߕ\vW�ҍ��IV�"�ہϒM��Y/�,��`��cݍ����7K�or�?�
��@Ҍ��ɡ���Tfܟ����"�E�\��"[����T|,���YP>}/��b�z>�����~�C�%�n�J�C���fS/S��iZ���a��2zܥ�aL�k9T�X��(�x���_�0`{l�k|R/���{,3n��P7#y2:ܳ��Y����ك"����I@���g��"�۟
���'���iX�Ȥj�Qғ���Y�3�/��iX_*�Y�$Q,��	,�X�R@��W�yRK#.�@��I�*�uX�� g_�_�����yX@����vV3�򰁝��.�ԜԜї˄e�2��q�gp��As}����BD�ND�ND�ND�O�g�Ϲ�s>�}����2��9���9���9���9������?�����B4�sN4�sO�7\k�K�K�+�+�+�+�7�a���o�i��E��M�-4Zh�ͅ�6l,�Y��af��/<���/<���/<���/<���U��V:�uX��c��Fx���<tg���ў:3�Fx���<tg���ў:3�E��,4Xh��a��E��,4Xh��a��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��uF���7Tn��Q���r��^���<5V���Zf�ǅj]��^�U�vkL֘�K�K�˳ah��|��E�l,r�UV��UZ��.�.�.�.�q���g\n����3Uf�h�s��������9w9w9w9y�s��9y��Uq��uo�u���3�V��7�a@����i�i֫�i������Ȝ��̌�FuFuF�X�$Q�ʫ���%�k���`F��/ݖaݖaϤ�Y������Fѓ��'��A$Q�jY�A$�I4JM�F$�K:F������u���4��{7�r�v�Q�(Y����'r��Ɂ�M�_pݖaߕcҰj�;eX��?0mqW�#�^1
�� �h��.$��<�T��n�7�@��V<���6�팇����,*;)<�!}�ª��1���*�|�a�nD1�Ȯ>ZR?�#�Z�?�#����#��_Q�������Ki"��>.;)r㲗(Y#rq�6������o��
�j��䫏o��E��VK�JŻ�KyovN�+-ڝ�S+��r��ݍ�"B⌬i�o��)����vG�+n��9eʒ��=Zn��/���~Me�ς[{ uir*�o�[��/ד�⳵�a|C����}][
<Vv�03m�����
ȸ�\vW�ձ�ݓ�۳�@챈k�vI��Aa��I�l�v����=cs?>6�c��mb�hY�r���ǊK�5Ϻ�jU.s�>)}-)#�R�.�Z�I�ek)C�d�9L�N�Y�S�V&+C��jr5kg(Yqݿ�V�&Ǖ߰�i��Br������4ʝr�W�i}���섅iyհ�r�sύ�Ɂ׷>����GG]�>x�L�2�K����I������d�4�	g��H���d"E|�	������"������3�����NO��NO���������������������ꌁD�D�A\ �W.h.h.h.h.h.h.h.h.h.h.h.h.h.h.h.hNs��8Ns��8Ns��8Ns��?��?�����C���Ӂ�8Ӂ�>��q�-.-.0�0�0�0�0�q���7�a�E��M�-4Zh��i��6l,�Y��af�ͅ�4��K�4��K�4��K�4��K�V:�uX��c��U���<tg���ў:3�Fx���<tg���ў:3�Fx��,4Xh��a��E��,4Xh��a��E���Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV����7Tn��Q��uF�^���9{�/|��c�ǅ��u�v�5Xj�K��f��i��5�<s���4N�5��9�<�UV�����af��i��d��s��~y��9��u�х�ӝ��7\�<����p9��p9��p9��������>r��U�^}mO�7����p�/��?��s!1�3#`o��F2���v>n�@�����7�7�O��c~��_s���'nɯ�U�UܓߥI97Մ
��1�aG"���F�{�_rΎ��d�{�)�ȧ�g��ڲ��z!ņ�/۫=�'���8���n�umۗ������ȻX�ҌY�v�Z�qs�_��9n⛹����/�G�L�Y�{�e.�zhVgk���®�/�)�iR��t�J���l�(zȘ��6����)Y/5�Dd�*��d[��y��o7�-��ݽ�{���nG�{��d�d��v��j�6�q#qH�n|��������╛�)Y�g�L�ɜd�dvO���G�&!�H������n)Z�!d���r���F�8VZG�$���?�D+ZnR��Y̷��p��5��D���Dɨ�?�.x�C�+��ۑj����؍�ogZΛn�*��ù`����`�p��ݯ�l���e}��e�nEW��_��_�7e})5��O�N��m�<:T��7)g�V�C÷��'�W�u�����k�!f)\��{��zc��b�ǋy��~*\tk��!�uN�\Eb�Z�Gkl��u�=FC�Em�*��K�[�t�f�yA��k25F�J�|���R�Pߕ7wQ!o��Jw+o�Y`�J[��6��V#��H��l%�����yzv�&�m��nR|;�u�oձ��g���Uq*�j�Q�Z�F5�y2:�X���dXݕR_&���g��dWᯂ�����6^OF�&^EI��3L�z�>��I4�h�ɠ��A$���D�'���$�RxD��O��,<�<� ga�I:O*H�yF�F�� Q�(�OTOTOTM�&�p��D�"n7��44444444'9�s�'9�s�'9�s�'9�s����?�����C��i��i��\n����WWWWo��}��0ߢ�E��M�-4Zh��i�6l,�Y��af�ͅ�^y��^y��^y��^y�玫V:�uX��c��U���ў:3�Fx���<tg���ў:3�Fx���<tg��,4Xh��a��E��,4Xh��a��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EF���7Tn��Q��u/|��z34ff��i����+XV��aZ��i�Fg=��^w��>��и�>��ם�y�kM�1��\hu�^s���� g	8H�@��W���g]�<�n���B@�3����|g��?����7c<���C�������i����'�2�q�g��p��DёF��>�'�H�n��Q�DݓA_,�W�+�����
<��w0.�Y߹g}�E&L
<�+����F�PK8���{�+��k�%�ݑO?&E�;���_ß>�+�5n�ʜ�.��v��c�U�Sxjӹ.�xj�6�ܧm�S����Ѡd1{��Rƽ���B��mܣXݻ)~s��Ѳܰ�\R����[���h�*�[�F����q6�6�K�M����l����-���<��?c����k>�5��-�������i){:���Y��ȷ��6�#y���kr1\��q���l�YΣw��\�v�^��dI|�d���I|N�s���q7)Y�ە��Y���I/��gJ�+���P�Y�J�"�e���Eǎ�
ԕ��V���k��`�	�����R�*�la���o�ܥ]؅%+M����q
�K_8��z��k+�\[���)+s�#~�@��H��K'�߂�j�`K�p��w��?��߯E�4v���@��`�����+?4���8-�4o��˷��'����I����<���_y�T:������g�I�ҶZ��t/����b��*\�C�t:Káߨ�����-ը�*���|h��y��aԨ����ң��+��������[Io�ps�_��x1J�
�o=��Kl���O/R����'N��E��I_�[�H\_��yU��F>5��e�=�*7)<�$�x���Ƶl[�����Jūc~�$�)��w$ַe�eT�l|��e�%��>���ѓFڌ�K#/�F��n��NE|�1,�I���$�%,�K"R�$�%,�K �xD�'���a	;�I�}F��|� Q�Q�Q�ѾQ�Q=Q7��M�&�p��D� ����������������9���9���9���9��������C����� sN4�sN4��uƸ����¸¸¸¸�}��0�q���-4Zh��i��E��L�Y��af�ͅ�6l,���/<���/<���/<���/<uX��c��U��V:�tg���ў:3�Fx���<tg���ў:3�Fx���<4Xh��a��E��,4Xh��a��E��*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*7Tn��Q��uF���{�/|���F���O66;Lv���cc���k�lnz'���Z?�h��v����ל�n/����<�.4:���z��F�_��a g���݂�|��_����H������H�7��8/�`��cv�&���bo����&���17~�A@�?��n��]g���*HE���e��k�c������_>Ok���$�U�r$�eU�p,o����5"�J�Ri�`]�d]����o����o�7��ܖ3��-�;��j��N�f��vʯ�8r��C�I�P5P�[�Y
B����J��ۆ��9~���r�?�����Y�[z"�`)۔d.2���r�.�%�WM�W�w;�w������B�{j�)Z���֩�jy[�f[��M����r��t֪8�1Mg;���e�=���k>ԹQ0}�eKicK����9{*�wt��F��g*�os��܎6���I|��s�φ;�2?/�\e�+��eq���r���^�%���_/���\��Ol����?@�=�c/�j"�Ƕ!��!P�� ��Jl���%e2A��4���V1Z�6K����$���uߝ�laPV�q#Sa��bGI�R���14�]�b��n�Qm�ek�-�5m�?�w�?���a��]�k+����yn+gw����yn-f�����.�
l�(ve�|R��m�6�C̥Ã��ȧqY�J���l*+��쩵��6/���r{Om��w���x4��K�p�)�h5?�R=���̇-��ݵ��?����V�d�]���՜�N�#@#���k/Q�od��wgL��w��ts���8YR�.u��=L�����yQ���\��t�N��E;�^�(��Wύ��+�n����+R���e�(���_���%,��6M �K�}V2(򡱺�d���۟V�H�[t����ݰj�5��)Tg���`�ݯ�}ư������`X߁c~���,o�F��)<M�F$щ4bM�F$щ4bY�}����g_:�)��N�
q�Q�Q�ѿԐ�HE$"�q=Q7��M�&�p��D�"n7��M�&�p��D�!9���9���9���9��������C����� sN4�sN4��uƸ����¸¸¸¸�}��0�q���-4Zh��i��E��L�Y��af�ͅ�6l,���/<���/<���/<���/<uX��c��U��V:�tg���ў:3�Fx���<tg���ў:3�Fx���<4Xh��a��E��,4Xh��a��E��*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*7Tn��Q��uF���{�/|����_�[�w��͍�Fg=�i����,����G�������~nn�3����J?�� g���_��}�/cj�2���0�c ���F'�����}���pP��K��W�}�v�6�="OH��$���o���'��7������o��|o������Rx�Ȭo����aw��4bO�R2%�u���ʬg�'��&��,�"�������t����'�"�쉻f��m��\8�6���
�p��rL�I��³��ʜ��S�T��v�;r�+I�G��{�|��Wi۵k�b��n��um�J��L^�Z�b˹W�e��~\[uo�nQ��U��N�����"�Ē�'�����U�B��Cn�kw����³ ��f��Y��X�WEqC��e�ǲ�hzj�=5X���?�q �u�jzǳ�7=Oߍdϕ�ʱ��I�[Ii�����9,>������l��7�gwp}ތ��Ky���|�a�Gd1���z7?^���w�����-�׷����{����ol��P$v_����$v_�K��8	"�%�1}�ˆ��D3�L~GVc�H��̜_����dh�q�Y�F���Kl,�+|�m�r�H����k���dh�)Z����W�{���b��C�#V8��)Z��|���t�>B��v��;����j_+nsO��zn݌*Eo�V�+<��+l�l�rj��[:9Y%��:����nr�ݨ�ë��u����U��F�ä8�.C�A���=�#��>:����+�!�[|>�-�-��2�S�|��?mO/���{��gv����}�T����||��T�s����.䎹�����h=k��e�8���Vz�S�#�}8c/$���a)�2߿���#��/@�i�\R�(R���l���~���N��$=f���ݫo�n|�)6K�����R��!qs�jĮR�6�	�Hȉn�.ʢR��%�Hϯ��_w>��}}܋�iq�K5���`F�#X��bM94L��3�D�O9<L��3���7�7�6I�I�c��XAN2�q�g�q�g�q�g�q7��M�&�p��D�"n��	�p��	�p��	�p��	��?�����C����9��p9��}q��\Z\Z\a\a\a\a\a���o��~�M�-4Zh��i��E�l,�Y��af�ͅ�6iy旞iy旞iy旞iy旞:�uX��c��U��V:3�Fx���<tg���ў:3�Fx���<tg���ў,4Xh��a��E��,4Xh��a��E��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV���7Tn��Q��uF�Խ�r��^�����̿[��33cf��w�͍����,����W��x/�`��	������ϴ~����a.��U������_I�Mc�2�t�W��ݱ��I|o��B#!��߳���$�17�FQ���_��I�RxԞ1'�I�xŇԞ&r����7�}X}W�NYvY�F�k�ϓUϓU���5,�Yƴ���ɮ�W�lY�y�ȯϓ�>O=)e��*;�+��+��)���������p�9$NI�
�B���Y�,����[����T�j��n������v��{��uo���Mܗ��f�ܭ[ugX�Swg�-����1|�����.ML�ҷI�SnR���U�����7�.E�]��Oc@����iohE6��(a��ui��������S��P�2UX�[SM/C�Q�ge⚛P�g8+�{-ql�u�g|ǳ�b�߶�4{;��ǳ�1��g� ���6Rm��粯��){Id1����piz�V�g*�kr8�܎6�#y���oua����[�R�g�v;���y���ww�/#��;ar�5��?�r�d�����o;�r?/��e#�;'@�v��÷9�B�\Oo�a�\e��v'�G����6���b�.YO��9x��Z�H��~K�(uj���p�-�;M�rt�m�-�q��I}�+����e;��V1L�_���9]Y[�b��Υ��W0����)��A�-��gK��uw'#~��!�+[<F��*����T�d;$R�1Z�+o�Hv�=F���=�Z��ju��v;s�S*yI[�l#��l�����
�_{]�bm��WćY��9^ܾ�eG�����+'�Z���b@Dz.���P3���L��u��)\�ob2:�d�՟�Ke�r��w*[9O���9̍��2Ҷ)����t�!HՏ��NG8��R�Q�ǥ)[�T���\������5���]�j�>\���We�Z�Eࢾ��ޭ����杯�J�ۓ�R��X�K�we{V�*�`�%T�U#��H��H�*D��g�F$�3���O9<bO���7�3�7��c��RAN�
��gY���gY�u�gY�u�gY��D�D�D�D�D�D�}�Bs�'9�s�'9�s�'9�s�'9�����C�����?�i��i��?8�q�m m m p�0�0�0�q���7��~�7��~�7��i��E��L�Y�3Zs�������6iy旞iy旞iy旞iy��U��V:�uX��c�<tg���ў:3�Fx���<tg���ў:3�Fx����E��,4Xh��a��E��,4Xh��U��EV��Z*�Uh��U��EV��Z*�Uh��U��EV��Z*�Uh��Q��uF���7Tn��K�9{�/|��LN?�p��V�^���݄�V
��z�<�֚1�4>����^

�LM�؛��7i#(�FQ���IF�2�e�˶�l#.�F]���'��_v�
���>�a;�����)�D� �_:����3�RNY�F%�)<Y�D�щjE��`������vUIFUIG"��E�܋�7r,n�X�Ұ�"������>��^Փ�^Y~����5��5��5��k�d��ɯݓ_�"��z�z�d��,mȜ�m������D0g�D%Jz������?؏�-���gα�:�/����Knz���n$���V��۹��"�|+���vH;����~*1}�uM�J&����l+�iӑ�s�H7mعyR�J�c��mEe
5B�FP�Q���e+�Ju���We$W%:�J�VJ���V��]<��G�+%s��n*9_5D%C�D�3���l{-�F�5��U$;�a�X\�R˟*YR�YԶV{]��cgK��mu�<m쫍��R���^�UK���vz�m���gr�l�^�n�q�W.*��r�=�u��~��o��]���l��B�~�#����ö����}�vÓݗ��j8}�M��y�߆6�Ƣ!e��+���H�M��$��K�7�O����{���������{l���}�ݽ��Wݳ��wwxu�-��)G��~�uJKp8�{�\���ꕽ���9+�,�b��ԏ��(1�g��镼|����/���=K��@$w�π�C)+=8�q+w�j� �J��w�O�E1:���{$l�U���ݽ�V��)#)���i_;t?)��d�T���g4��w)��9&��x�o��C1b�zYY���]k���v�?_cd���+Y�W8���������}��vO�#��>����������d�Wi(�����/��� �WBG쫘t���::��Wk*]�W�XO�S�����������T�/"H{,�Cu��͓�+����&"\�T��:�^�	�`Ȱv��A\,��e#"YFM�A$�4baX9��-sF��XD��@��4s��$�mZF�Z��a��Ff}̓Af�����M��v0���F�Ay}�Bu����~y��9��?<��������i��i���w���w��|&4&7�O��s>柜o6���ی7��~�7��v����͆�֙�4ch��.х�
�
�
�
�]q.�U�]�]�]�]�]�]�]�]�]�]�]�]�]�]�]j��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��UV��Z*�Uh��U��EV��Z*�Uh��U��E�^�2��՜�Yբ�EV��Z*�Uh��U��EV���Y�՜�Y�՜LN8(+_�����>h��/	��_=n��>y�s<�'[�_��AQ���2&q�3���62����#n��N�2v1�����d�c'_:����o��]��}���a�a�a�_:�)��+��x���g,��Y}�$�Q�4bY�A$PI�%���J���Dl�#g�I~}%�V7t�n�X�ұ��cwJ��V�R2)�*���z�y��/זOV��'k���wd�}�gd�{�)�W�d��c�D�o�O����'�����!�8�Ფ7!@�[wQ}�7u�E�Q�)�2(���i"辪/���!��ob��:��x(V�8V�o��Yjt�i��v����U��7m%p�ߍ�5�jj�MV�*B�����(U��R��J^���Q�ݨ���
����J�I]�-�[���J�w%Vߒ�]��Ed�qY+�vJ�]���r�5<���"���C�D��V�L�S	�D�9Q�MdlYc�I���<?Y'��I�\�eK�_�Զ2�>�M�ɪ[94g�����y�]��g����o6w-��wy���ow}���v��wv���M����p��������|�\o��k�����*^�˞�r�ݹ�w ��M����D?X�Y���o����{r����|��Ɋbh���ϕ�A������Y����v���$>X��]>��o*~��+9��?�p<ukQ���rX@���y���jTtS��`��Ih�)�`�j�T�s���^ץ��p0��s��v��Ys���C����"Y��v�����v�M�*���V~[#'���݆Ι��{t����2:��r�)���E�P���s�+}����ԭ�?a��<0}��������vӡ����鬒��T������b}P~�و�ä�j���Z�$1%t�Rr�M��҇z��x`�g~w9��A��ܬ��a��Es ��1N�)y�J�\l�;{*�ӴTe����d8��Q����n���������k�=yo��a��.L�MZ���U~#>�ÑGVN�I��uW�5���!�%Y<M.h,�oTO��ȿ��I��Җ@���,����4&�'7ۄTL
&��y�?<����s��~y��9�����C�����?��w���w��|&4&7�O��s>�y�����0�Zh�~l7mKյ��7sa�5�kM٭3Zs��i��\.xY��af�ͅ�6l,�X���������������֪�UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UUh��U��EV��Z*�Uh��U��EV��Z*�Xe��/|�Y�՝Z*�Uh��U��EV��Z*�Uh��K՜�Y�՜�Y��ႂ��������		G�%/�b`���Q����77H��|��?g�t�S���$� �c}�M�񓯌�|d��'_:����o���_:�)��N������	_���O9<bY�F���:I��NM�D��)dJ�%g��YĥQ�Tc"6y�ȍ�Dl��/Ϥ�>�y�3ϱ�}���g�c9U#"őbϰiW�d�Փ��ȱdX4�ڲv���&nȧ�f�8�K��o�*�$�}���eWv�'Ƀ��7h���C=�+]
�B�g��8�E�n��C�IϜC����D2)�;*�ʮ�I�´�d����eȦ��ݓ���w�<�B��~ﶷG' ђ$+�VU>BR�$�!-����+븻��]ج�|VB�+��W���YAo��A-�ԬZC�Ε(]��2ܥj[�1��,��*�vJ����\�rTG+惕���?��hyhf[��-�=���jbb�h���=���e�b�h��6����a�+v��紓�m$P����i*��iT���-�dc��iR�:����/c�����v;�}��/cŵ�ܶ�;��[ŵ��R����ogƷW�g�K�rT��+��s�g�R����z�mn��{����~����~�ը�p"�T���Ϡ�r(2��)%Y������+���p�^@x���}��G��Y<Pc�!eq���X�v�������<���d��Y��E��>!�^F��u{��-�=��-�w��cn�l�T�t�Z�d�t�^+��K~��+[��6�)g����g�c$ku����۱��2��"���wu��*�&���ǣ ��/��>r׃�x>�x����T��5?�K�|�^����|�|m��lz|m����\����ϧ���p}�s�w��^+���]
^/���{YC���t���G�|5+/����b�x6�S�5�Z#+6x�'V�����qt�
�d��r;[�d�FG�_����||C����bwj��}�q�õ*n�����Q�b%���қo��H\��$�ֽ�V1��gw�>���d��O<��"'�'��$�>g���Y��}���p��F\#z�:э�F���'9�s�'4'4'4'7���t>�}�������Ӂ�8���~q��@�@�@�@�u���3F6�m���͆�l7sa�j���_j���1�c�ǅ���������6l,�Y��af�ͅ�]�]�]�]�]�]�]�]j��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��UV��UZ��Uj��U��U/.��K˥����yt��^]�^�2��՜�Yբ�EV��Z*�Uh��U��EV���Y�՜�Y�՜LN()x()�j��W�ڰ_j�}�j2'�J?��	?�P�3��}�����F�F�F�F�X��c}|d��'_:����N�2rx���7��N�
u�S���������O9<L呩djMI95$�ԓ���Βr(Ԛ1,�K"Vq,ŜJ�%��F%Q����F�"6y����_�c<����>�y�3ϱ���*�dX��U�*����'dX2,�v���"q`N�~ܪ����'�*�$�{���_��w�>���0(��Q�����v�*����~i8t�:M��l���0(�`Q��rJ�Ãm��$�3��*o�_�*�հD3��$-]en��V*b��^ֲw�N���V����>P�n�.ҥ+�<\�����s��$�!%�,�9]�λe�vBWd%vBKx���R��B[�$w��S�HWm�ZT�������Ue��[~K�%����]�h��\�W:�#�O����Q�\Ps�hy�4=4%�MC�}�i���h(�v&)���k#b����6���r� )d�&�r�a�����>��թl��[,���>��Ճ���-�WeKe��nA���}��Ki�R���m4���~�J�ݹ�w ��ږ������`���w=e�c�s�`ǳ�pf��a���)Կmٖ���3���)����#���|���0b��C�~r���B�tR)���$���/������ʬ#4N.V�Q���yJ�:�ƥS�v��)��|�!��qXb�Q�"�:��]�I�uf�C���/�����~��+[��6;L��M��jq;�'-��b$-�vP��yY9aO��ry*�6�����NK9f�%��伎��^_����K$�%�/��)"VǷ����W��ΝK;���{]ON�������7N���q�^�D��|J:��Ѓ�]�Х��0y��pw�����/|R?����{�BQ�I]4��"���ކ4�8<���a��w�R�zu)���x;Y��zm�Lz?����8�����P�v������P��G�l���n/)!{$~�Q��ՄS���HR�vn	���55�<��##�P�c�ө;���}����l#(��]��걄��$��|�I}'Z1��������������nn7���o��ZZ\�\�\�y��@�i��\ny��1�4N�C�g<�y�1�ch�ц��o͆��o͆�V��j�V�Æxp���<2�ᗿZ8e��/<�Y��af�ͅ�6l,�Y��af�ͅ�6��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��UZ��Uj��U��UV��T��^]/.��K˥����yv{���/Vr�gV��Z*�Uh��U��EV��Z*�R�g/Vr�g/VpQ5`�j�DՂ��V

�߷~���22^6
�L%�/���8H$
'�'�'�2I�I�c�c�a;)��+���J�%|�	'���&u�J�%|�����	,�K#R�Ԛ�rjIɬR+	Ȭ'�c}�$�Q�4bM�F0#��%g��J��Ī1�<�FE#"��HȱdX�,Y)U#"őbϰiW�d�Y;^Y=);VLב7p,�2(��Q�իr�N�*�$�|����7������'�gw{��`_���ې�9%K�B�*������ɮ�I��Ȯ�Yѹ`U�H��K�g���!Y�w�Ӌ�c��dZ��n��ݲ�(m�Eb�E6��!K֥,1�J�*P�!��-��e%vREqj섷�R�!�R����eHvT�!-��!-��!)��!)�U>A�v�}>�F;e��)_-���*6�B���ߋ�]�-We)z�/���,59*�G+����A��T�#�;	A��P��m��(��&=���r�(z��Z6٩���d�=L�٩��jpcڜ~�J�҇�4���[��^����n|r�*[-ږ�w�e��׹��{,�v�"�ϖ�Rʞ��ȇl��z�ZM ��!�i<W���������ռ��0��B�m�����w��5=:�E$�����}���c��=��+�?9�}�����6���?ldWg��_��*��kt�*��)J��m���vH�Ht�����bq5o�����{�m+[��lv��oʻ��۶[*f�SY�i�:l�^J�we^�B��r�R��
�+%M�el�,����ew�T����yQ����e�)�nJ�!B�`�P$��,��,,�W?�VP��{���QL�N)z�Y^/+ީd�79C�s�<0|����� �����Ӄ�^���ӽ��WO���x|�S��A�������t�+��ë4�-o%.���ӡ{d+��� �z�B�H4-��Yc��
Q�b�{Zܯ�j`ſ���ܼs�!A��G��pqNU��
�m7��<�;g�����d9#S�]��{�kz�/!�>u�w������v�YT��$�Ko�'�o�o�'�$�`o���I/I/������/�q����_����	�	�p��A\ �W+�����>x��Zf���z'�3�g\ˌk�k�k�M�-4Zh��i��5��Wڵ}�7ma�/�����j��w6�Zh��i��E��M���af�ͅ�6l,�V��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UR�R�R�R�R�R�R�R�R�R�R�R�R�R�R�R��2�ᗾ^���έZ*�Uh��U��EV��Z*�Uh���^����^��>��F
&�MX���PTa!/��q15bbj�}���L%�/���?�g����RX�N�����
vS��W�+���J�%|O9<L����J�%�Մ�	&����rjIɩ'"����r+	��߃aw��jM�F$ь�bE�A,�Vq,��1*�J���FE#"��bȱdX�,Y��}�J��'k�'�,�d�}�)��70g�*�nUw�"��}^Z�X.,�o����m��\R'�|�n��
�v��[�-��r�r�_�&���|Rk�$��Ȩ�Y�۳��"����[ug�Yw*Ӵ���e�p�M�C�~�̃�' ё��kX���]�t�v�(N�!)R�)+��+�Eqj섖�iʐ�A[��ʷYV�	n���	n���	O���	O���*� εe�j�;t�9PHx��<]��vC�Ր�+��vC��-�e�B�R�]��범�VR�o��T�jx�5<G����;	C�}���r�5=7ڞ"
+����j9�=GM,��d�4�=�ȏe���l���J�׊e���������k5a��X~�J�χk%QMd�=����$�̶SY*�e�U9*�+(FP����8�p�j���l��&��[\���S�86�|z�-���_��pqJ��VP}\/����/%���C��c��G*Ϭ6Ma�Ku������JEI����:T�o�e彆������]��ݐ�����eL��mf�)��[�^�~'Q�|���Ο��H�m6'%l%)C[!Yv�YK{����l��e���u���+'���6Y݆ӕ����+T~���ʕ?�Ij���)g8�K��=q+:?9�z9Y%�r>����<���E3��d��J�K���a��|z�܇S����/ ���Jw�)[�äM��Տ/�D:w8or=�\��}5;�N��ԫ�й��;Zo���C����;�s��_�FN�����d���x��R��Px����iq�T�@p�^֝�1~�tC�ƶ���N)����N�V����5����~���&�~��%'�Ht����\k%<�ܩb2��n������+8�kJ�r�(�hΨި�o��y�c�^�����������/�q����>�!9�9�9�9�9�9�9�9��@�@�Ɖ��=��6���5��Ϟg\hhhhk�k�M�1�Zh��i��6�a�6�a�k�Xnڵ~kM�-4Zh��i��E�l,�Y��af�ͅ�6��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��T��������L6�m0�a��i���{���/Vr�gV��Z*�Uh��U��EV��Z*�R�g/Vr�g/V�� �|LMؘ��~����((D"'�� ����'��!��O�O�O�I��N�u�o��}|��_:�)�>�Y�r�$�	'���&u�*��|J�	a��I�Rk��r+	Ȭ'g_}�}�u���]�RQ�FݖF_&���2�e�q�dPIE����L��g�~c"��HȱdX�,Y,�E�J��^Փ�d�yd�$���߻g~�����x�h�`�����*��*��fܳnY�dN)���"qH����r�9%���D�rY�,�R&쉻"��r�9%��c^Y=Y�Vtxp(�0g�$ĥrb7��~Q���������镊��jC����O��O���U>BR�$���vRKx���Kr[���\�<\�<\�<\�R;�R�$w����Z;�Gqh�-ũ��!+VT� ��$H(�-ũ�U>ʧ�3��3�SU�j�eS�$w�b�HWiX�2.ԇ��-�\�R�9%q-�]m�W�|�滕�]��%��$�%A[�5ܬm�ao���qz�"Y��Ed�UO+�S��Pd���#J��Ҩ�4���Z�J��ϡ�TFM"��T4�=���r�b��:�V�+���e�߯n�Z�J�^@�:֜�����ը��b���}�Y�Qg����b�)��^K���}+���(v�� ����kL�V�(�p65h�ynH�/K��Px�4>Y�����l���X�����D;�ݐ�z���$G���ef�C�S"�Z� ��*� �g5�1o��d;uJ;Z��2�:�N���ֲ�*U3Q���9nH�Ht��F�֫5:����s�##.�<�H~�f��S��[店�A�[�������L����I�s�W54���}����������B�J�)�E-�������迪=����ߐ;���P��0�]�/ЇP=w8�����C��J78�
[����J]:Z���0�oN��"u����qyj��\\������W�s�Y$|��P"5�6##����+�Hw*����$1����e;5nT��wag�#Y�����lW��#��m�~N?����Ƿ���*ܩ���X�ùܯiW�lh�|��pP(.���8.���8.���8H�@�����/�q���n.��]��������?�i��>v���~l7y��^v���>��i����445�5�5ťŦ�m�-4Zh��i��66lm�-4Zh��i��E��M�-4Zh��i��E��KUV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��6�m0�a��i���L6�m0�a��i���L2�ᗾ^���έZ*�Uh��U��EV��Z*�Uh���^����^���?�AA_v

��g��	���
�q�W�A_�q��O�O�I��N���o��}��>�>�>�>���<"O�'����O:��|J�%a��XA$�)��V�XNξ�:������ݳ��"��&��,��M9e�(���nȠ�($�	g;8����2��Dl�),�E�"őbȱj�ڲv��z���I�ݑ]ݳ�rΎ��:;�+��+��+��+��+��w�ȧ�"��}�f䱻'n�۲v���'qI�R�$��,oɛr'�{�)�ɯ�OrX⓶��)c^Lݳo�(�c!e�enMO�N��[j���Km�bu][fV�Um-���O��U�>��YRܡ}w%FC���T�!)RC��!��-�ҥ+�҄�҄�҄�҄�҄�҄�҄�҄㸴w����	Z��VT� ��*�!)��eV�j��+i"��+jԂ�YT�	O���[��[u�^�!a��X��8�/5�P�J�.)X���!��<��R���Q6�*�[��%�*�ߕ���d��g!�ܥ�o��k�)Uw%*��Uܔ�+%dWrR��K�%Y�rRh��'��Rx�V�[���eȬ�S��a��gL��o5�4�t^>�,B̈́-㻺~)��8����P��J�_c��j>r>+ܑ���%�^5F�#�p�:G��g�Q۹�c�܌����mk��w���ŝ}��f^���덯s�g<j� �I}���!���R�*u?t�!��qXb�*U.���]�Kt�=*;�Z�#�I���Ku���J���pz�*S�C�4�}�R�V�ގ썿��	{�]�[5j�H�3»���0�8����C����>/��//%��[��]�qO��n��ӽ�?�^���B���dR�#�Ȥ_�A�{(��+��z���{~�~xa𯝳��l��C��|7� �@t>F��|G娤BQ�P#��ls�?�B�0���-mi��n#���v���.�d�S}^��+�_T;�@b�+'���P%b�-{�J?+���ݒ�Ԥ6��ﲽ��KkOۈX�vREB�l�c8�G�+���Ͽ�{m����!�Q�\싕���*b8tYv��{*ܥSϯW�# _t,|�����`V0(�d
2���W����_qv�������>�}���}mO���0ߛ�v���W�<�]�j��/��8��������q��u����g\�y��9�<s�|�Ϟ9��>x��E��M�-4Zh��ij��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��U���L6�m0�a��i���L6�m0�a��i�^�2��՜�Yբ�EV��Z*�Uh��U��EV���Y�՜�Y�՟�/>_������AB ���D�D�D�D�D�D�R�������}'�'����������"�'�I�ϳ�}��6�2�<b�%_��%��5$�V�XNEa9��V�XNEa9���3���O9<L��3���M94L��R�$�	,�Y���&vq3��J�/�X�Uc9U��V3�X�U`�X%V��D��,iI��"�VE~��܊�E{J��^Փ�VO=Y<���I�ד�k��,�}�J��^ү`�;$��H����Ru�XձvX5l��=�)�K6���&mɝ���P�e�o��.�m�u��4۹:�����"�v� ѷ�R5O���
� �R
� ��
�e[��}��Q�
r.��:�5Z�V�]��J�*R��)_��O��n��J�.�r�o%V�(]��S�YT�j�MS�%�P����vRj-�T�G)[e+iR�������J�)[S)�ՕO���b��X�T�^l�n�2�/Z�q�d-�
��!\Gl�c�jA��H?�R�|���e����)R���)I�z�x��V[���<^*B���x6�K"��ϐ�vv�,�; ��X�<W%&��RynP��Y~�e(*����c�8>V-��ޑ��j����wv#��tY�Ӗ���?�Ju�"S�1*�;��k~r>���$|���9��,1��|xYP$~+�|�_~�K��s����ļ�W|2�=%��X�vF��	Uw���rE��z6q�O�+��K~�D���H��mj�O����[u?�C�A�ۜ�!��T��S)��k��m�Y���R��e���5�=��'��e�9-�"B�IR*R�yYmw;���B}��8t���ҽ��I��lC�U��'������x<G��+������a��Q�p2�V[�rZ��Px}PT��[8}�>�-o�zj<=}���W4��e��C��P�����{�����ߞ�+��w�\!�D%Q�P%��w��x�C���s���-��oz��T����R��jP�j���yj��v�	ky��D;�X�������k����PL&KI]�ȵ�=�A��t��R�Ѐp���5c�s���eq���:;�A��[�_d|v+(vZ�_s�[�����W�il$�r�gՑݰFZW�k����`�Ձ���̸¤�����8<�]}��i�]	��N��K�熏<4tKݵuj�����ם���s����H0�8y�9w�wa.(���i����3�f�M�-3af�ͅ�]�E�<s��}�k�㞋L�Xh��a��Uj��V9y㗝��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��T���������kXֱ�cZƵ�k�6{���/Vr�gV��Z*�Tn��K՞{�a��^�2��՜�Y�՜�Y�՟�/>^|�����AB ���D�D�D�D�D�D�R�������}'�'����������"�'�I�ϳ�}��6�2�<b�%_��%��5$�V�XNEa9��V�XNEa9�����J�%|�	_�A%�I?Բ	,�K �q3����L�#/�R_*����r�ʬg*����r���*�J�v|��&���zR��V3�X�>����X_�a~�}�Z���7��5l�z���ϲO~����Q�F}�J��&����[���v����.�ƴ�\�%c]!n��&����>Q�&�9�<���JUd�B^H���Sn�+s��)BKx��XI�j�����j� ��U>A�2��+i"��+j�5O��ػ�9J�N�����F�)��jAS��:Ԃ�H*|�����Bv�A!��--�W�,�~W2��S��j�mS�+�1�N���U�³XVm��}����Ֆ�>˚;!h��y�l���޴�oZT�J�"m�M+n�#d<���%XWq�en7)M��Sd��,������	P���
�n�+��[3�4�[��c��Iol�X�ڝ�Ɋ���T���-�2жVb"̗�T,��?��NM�A�k�����]q��W�(^��F�r��,� ��u�=��,�n�+�i��.����^5��\�e����*t̝�LmO�)n�P�;	oۭ����~'Q��iRT���b=��MF�J�[�����G�U�t�$@2y:�a�l"�ߕ+[��2X��#%��b6L�g�����}���Vu�9#-����qE]��`����&��kQ%�2�/�W%��$w߲i��X��;��w:~.;8�j2E�Q(H��+��>[�㲒�;���}�mO��A�ԭ�>H��ҷzp
����v�4O�l���8}V��U�����ǿ;�HWz)
���	j)���\!ЇC}P�oN���~�>/����>"���_�s���(��@�jP�F�@�A�ͬ*Z��K[���)��FX��[`ڟ$�JY�_����٫$�ޜ:�-A�d�b��m�:��ߥөG���L��)���:�#�ږ�"ݝ����܌�Z�wrVTq{*9Cu����u���?$IT"7
�"���gܰy���}����,ȝI����EWۋ��u�8���<��U/{�9:-h�=�U/U�36[��X�٥�q��:/��хq�q���f�M�-3af�ͅ�]�E�<s��}�k�㞋L�Xh��a��Uj�������UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV�����������<�ǚx�Oi��<y��4��߆^�z���:�Uh��U��uV�^����k�2�ᗾ^����^����^���y���������3��|��|�'��|�'��|�'��|�'��|�'��|�'��|�7��|�|�?�?���>�>��_9de�����3��W�$�3�F���5$�ԓ�RNMI95�Mb�X��+%�������������O�,�K ��$�&rh����2�U%�K�T�ʩ/�R_*����r��F�lX6,��*�dW�+���m�����UI~}%����F�>�z�7�W�ݓ�ݓ�쯣�'��_�����U���R�Ԫ%*�\���)>��;�.���~L�ʕ�
�vP�*P�!�Tk�*5ܕ%v������׶?�/wam���_��2��>���umn�����[I�2�:T���e����js)Ne)����V�J�t�|�)Q��Ue�J^[���J^C�*ۤ�r�ج�V���C�a������R;�V��o%VF�$kjC�0֩���v.�T�vC�]��*4�]t�V�M�L�_L�_L�_L�Q�)��Ec�XÔ�摣�����o�"��H���H?��v.
;���Yi#�}*P�Kr��C�%��-��[��[`����+)X[��R4_D�@����\N䭡Ӣ���8�G,r��[�r���7O�+
Vb����<jl����2;��q0����e2���]���[ވ�?;'{�ރag/ �Ht��+>s≗��3��Ykd*%�5w�'Ŝ�?r:�J�l0$�o8����}��PሥFG�(2>�o������ʕ��Ku�����褬��$t�!�����*�R�S"��=�C�V�|v� �z-؝��$bju��F;Y��k5:VR�J�-����e��Ay��d��I���@ݰ��e󲏏�l�\�Y��)����V�qZ����\������"���m�W�����[]���[�w^V۷`�os�!��i[��~�]�W5ۗ�+������|�ʎ�/C߅�{�:·��o�c��;f�B=�Џp�#�>�*�D:p��t!��>Ї½p�W�
���878W�Q��J5/�F��(Իc�]�Gk��p�7�؎ַ(��*��>>�m�}+s�����"Y��z��>�s�����_��]J�܊vp`�~�����pޟ���~g�L�H�#^ʍ��$�R�(��/�&��!.}�;f�M���)��&�����"���nÊ� ܺ�wn%Q(�l
G�ig��gW��g�o���qi�]��޺0��/ϛ6g=��_�:5oK�y���^x��c����s�硣3�f�M�-3af�ͅ�]�E�<s�|�Ϟ9�ͅ����UV���������U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj�_
_
_
_
_
_
_
_i��<y��4��<�ǚx�O��e9z��EV��Z*7Uh��������/~{���^����^�����������?�g���PP((

��A@�|�'��|�'��|�7��|�|�?�?���>�>��_9de�x���+���J�$�&r�Բ5,�K#R�Բ5,�K)�Ռ�	a�a�a�a�a�a�'��A%�IdM94L��g�~m�����6x1����l�iq�8�k��H��`R0#Vq+8�����&x��Dl�#g�<�K��.�W�쯣�awJ�y�H�2�U��d�L
7)3^1�ߖ_��V4���Ԓ6VY���z#�T���H����InAGkjea�����fA�'M�$Je��m�-O��2���T�%F���-�g����md��o%�;!U�$jAGd)�x�۬�"A[�	�e	�d)��"��V5�Y���MGd�!%�ZC���*� �R�C��J�vAGi��KvR���֫j}5�Q�O��T�mH��2����byJ��eb��X�Z�f�)��w9"�֙m���JwZen� �֤�J�R��; ��r�l�(X��V5�J��(F��5�m�fV�m�񬰨�އ��8g�Ź�#�#�.�1[��tY�d���P�1!w����+N��JE=�n���VIT��e��s�얥o+aԪ���4�*����[:p������a}��R���GO��u�,�\�7��V�-��IX��[��b��moc(J�
B��]���;��۶Z�fӕ$lv5���H�e�r�����u�\��M���2�*mc-!SyRU�c%Yv9[.�J�yY[.�M��쳻�v��͍��v�-Gwicqvª��|rV[>=V�;o'���r�B����q�o�+}�[��=ح�g��o2��uj+e��/!����gGO��Ev�z�$J������{�̷�\�{������^����Q���n_:��A��;p���P�o���E9:qM��ӊo� =B�ހp�����~�������n|2�?�Q���{�؎���C�����!���P�;8����F?@�{�}{��R��\P�S������p:p~�?^�g�nw.�{v��t�]����n~��ȧ'z��k�.���������n��c�P�ݫP-�^�=6GV�5���*ǎ�� �治���V a�>���J��[ܗ��Z�����j��;�;��Db3]����07��a���/�

	v`h��v�5��-��q���Wn4]�qw�������3E��M���af��.ͅ�E�<s�z-3afµUj��U��r��/<�o͆�UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��|)|)|)|)|)|)|)|,y��4��<�ǚx�Oi��w��e9z��EV��Z*7Uh��������/~{���^����^�����W���P�3���$�����������:�3��:���`o����g���|�'��|�'��!��O�O�I��N�
vS���'���
vVU�I<L��3���O9<L��<bO��$�%�ՏՏՇՇՇՇՇ�|�g,�94�h+��Wȣ/���2���#/���1���YĬ�Vq+8ŜbE�D�Q)E�A,�Vq+8��5*�iX_�a~����3ϤdF�bXL��Y��kػlݲ��j!,E�l����o�it��C�\k ݬ�({r;)��!8����b���˯�{����R�BKx�z��ܝnտ;S�F���j�!_�λe�� ��ԑ[S)�e9��$j�)XI�*BT��9[�8���Z�!$�j�[S)�"��Sn۩�hy\t+NR�S�/���9IQ�����Tr��e%FJ�S�Q�쳷�W�rC��9	J��VU*AR��A�� �H���jH�����U���-�U���e��Sn)�޵��đ[�Z��Sy�l��^v�m�>��H���E��(i�|4�����N�l�y���/o���	^Vgey��d�J�ShP�:�$�+2P�GIT-���*?���A�/�Ʒz�b��z(�+�Qo��d��,��?Gl�۷,#e�Z���:�ʡx�?�a��I|^޼L�$��vS��7��J���Y��4K��;��ov;��e4�]D�!wrR��c��z=�ʕ��W~^�v�g�l"�=�?g���YL�Wa��{r�lN�S��gr�lG�e���vYOnε��ֱ=�|��S2��˕���e��lJ;��i����%�G/Q�G$|�(�;~Z�!m�Kq��K�ze9OƮd���H��In8�B�Y��m��?-��I}GK$v�1�HY#g�y<�`{"�.^���۴�lwJK[�k�V��[���z�m�^����^�^+���}�=�}G_�A��P{=V��U�r�nz�����=�ӊ\�qN.�z�ފqz�/\���m�a�|v������������Ƕ����>VH=:�l,�iz��އ����?���Sw�s��|n@p}Ϝ;_���T�z���A�9W���nz�۾���
���>t�r��ܶnt.|>����r����[��h^��|[}�[-q��~�8>ͬ�+�~v&��ϧ�$\6G���5Gѯ�������V�+��(�q3��y���3w���^&�����蛉}Xh�c�[�����-fh��i��E�l,�Y��˱˳ah��i��E�l,r�UV��������6�a�6�UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��U��UV������yt��^]/.��K˭Z�ի�Z�ի�Z�ի�Z�ի��߆^�z���:�Uh��U��uV�^����k�2�ᗾ^����^����^���?����	8H�@���������:�3��:��� g	8H$

��A@�!��O�O�I��N�
vS���_;�����$�&rx���g'���&rxĞ1'�I�gc�c�c�c�a�a�a�a�a�_9g��>�M|�
�4�(��q3����L��gg;8�����%g��YĤPIJM�A$�IE�A,�Vq+8Ī5*�j��үdR%T�TbU�F4�Rw��#��y����^�no�+�>B���7x�7�#�=�Y�9)'��\6����H0�8�ř �	Y[���FK�}����gQ�\[�p�Tn��'�����mPrTm�*��+{+j=���\E2�c����-���:}5$VD}Z�#��+�YT�ڙ[S���Xc��+�ϕ���l�����ʷ��YIS��<�+�Ht�Ƴ5�S��[��n���qò��̭�ISŪ8��)x�V�vAI)NVc��}#G�Km"���m��[e�1��8��^�N?v�m�L�Q�V%�Q�4�m�J�P����1Zm�/q��W1^،1(HS- $v"S�,���$����£�xoC�/��8�|7����ϻ����G��ޟ��l�+���`�O�r��NW�ۢ�IBBݰ���>W䛣�z%~:�܃�?pT���mژT���]��k�|?; �Z�V��8B_[��j=�w[n�죻U>J�l6�I#i��2�mF�S���m6'ѽ�HR�%��d�_,^/{(H[�*R�IY.졋��8���F�ld���H��r�-�����1:ܥg{���_7��������}��V���{a\��^���R�|��=��Y<NS��}>�C��=2^�+�Kt�f@T�����d�{J�8��W2�����>V<|�*�i�<|�*��WGO����T��dW6���*��z^�~G�ߑ��x���ʞ������*:�ʎ�΃�����}��g�����t훽��B=��nw��]8�z=r�E8�)&�
�@;{�8��)r�Tuc��ޜ:��P:{X�����t���;�g���vt����g������0�N�?���T���=.��N���ɽ6���އrw*:�K��C��E;=u.O�Ss�l��=�}*�����w}W?�^+����|4�����b��?��+��퍌��ix�^�����#��+�&��ݔ���)�hT�crO�J�%�����,�xV}]{�"Ú�v05n(������j2�{M�-4Zh�ͅ�69v9v9vl-�-3ac�c�Z��/<r��/<�o͆��o�j�UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��T��^]/.��K˥����yv3Æxp���<8g���{���/Vr�gV��Z*�Tn��K՞{�a��^�2��՜�Y�՜�Y�՟�s���/�q���:݂�v�߷������n/��|O;�y����H���$� g	��B@� Q���Dd"2�q�ga���������v?�0���)��o���|����J�%|�	_����� �a:�)��N�
u�S��������g&��M|�
�M�4�h+��Wɠ��A_&���&rh�ȣ/�F_&�I�Ȕ�	'�W�H�R(��b�1g��`R0)�y��0cX�֕{�Ώ�_���읗=%n-�W�v�O��g��c��\��o�+�����I�(�+�ߑ��m�9�6,p��b�/!@^:B�t�x�,�1LV�܀B�{g��/�S�;ȿz�
��<�1!���V���*��$=�Y!�����q��g9K9YL��5�-�8Z��Uݮ�7ƶ=����-Ky*�9*�S�y���r�-��'k���r�a�kQ�IS�YAR�U�eV�)��x2Z+���h����vROP#�nF��=0~V�v_�-kk������l� L�콾R�O�gZ��Z�ݭS�֫xd�t�2�W)X���]�V'L�_$S���4B�;M�y���5?v���(p�'A�d|�efJ�$���G ����/B��z����oW���xZwG��x�[��"�{��b�I~��G�d��oJ���i�:�mb&��n�P ��Б�9NGj>w<GCy���
����F�I��+a���vr�on�)T��s�{Z�Vj=�m�e��6��~_aS��h~�m���d�1]��C��i���+���D�n������"Z�@2x�����kk^��w�j;��Ι��H�-����d�^�"�L�����̑J��j�}�C�l����͟���x
�M
�@ݦ�;d������Z�{�9&��0�sO��N�{�	�����*K��/��ۻd�*�12iY���r�o)&��.�H�r�D���Y�j~��Ƞ��� ��o��m�>���+�����9���������*:�ʎ�r������{��慎��n@v��=��m�-�]��~����pnqχ�Q���;;�<��o�=��n����N��ܠ�g�)���{"�P�OW�Q���x��z�߃܊vz����~���*���7����n�#۾~ߊ+����qM�}W�S��îQͬ+�Aծd;?_�����\��}P/W#���vͿ+�\��=���|���Tx�e38�ʠ:\��gd�BO�`ۤrW�݌I[th,��3������qR55�}ZKQ�8Q���F������3љ��E��L�Y��ac�Z��.ͅ��E�l,r�UX��^x����ߛ�-]�j�UV��UZ��Uj��U��UV��UZ��Uj��U��UV��UZ��Uj��T�Y�՜�Y�՜�Y�՜�Y�՝Z*�Uh��U��EV��{���/Vr�gV��Z*�Tn��K՞{�a��^�2��՜�Y�՜�Y�՟�s���/�q���:݂�v�߷������n/��|M�'��n�3��B@�	��B@� Q���Dd"2�q�ga���������v?�0���)��o���|����J�%|�	_:�+��Wd�Wd�7ɠ��A_&���&r�dY�A$�3���_|�2�|�g,�9g��>�Y�r($�	�w2�ŜJE��$�R�D�	g��Yİ#X��#J��`ȍgƷ+Ь;��W��WYg��m����q��mk���P��J�\d��o����m����#���"�)�B�rP�_����~,g5�[#��c�tX�nZ��K\o��?�����e*���R��)T���^Z,��G��Ds�G���@{̯�y(B�8����r:B�g5�_Х�Ф�_O����)z�|����Ij/S�c�0J?��H1ԅ�$����[|5(�/ �A�)-�x���Y��5`/��ә-ݖ�p�+%:����+vp�gd��өv��]ȧ'���Х�v�.>+���l�~����r�b�h��v�٦���#hzhJw�;�)�����{�>���B���r��A���'�B�V%>5���Dj]��mk�(��{�������\�:WgK!�zi{IF�G��)�}=���.��G<6O����~���W��S�k���0]d��F#�+%�}/��b,��Ͻ��m�����S�� ���N�c%r�:ܝN[��FI�9LL�S���4{����u�\Thu�v�K��}Ժ_��5�"=���m�����#���Y�IzN��W<�&+���6<���c��z#�?m*����H����4W)�[�2�c�J��r�m6�I��s�t�݌�����-C�t��E����c�خq-t%yG��x{��O���Y�.��.Y��W����y�9�Ճ��g$ig�#I������K::d���$R��g+i�j敁\�vu̷"����v�?ݾ������^+��s�x�����t�z���������:�:�����vz�{��f窇r���%�f���ܮ��m�r�K�� ׈�\�;f����x���Ѐj�aھ���n����^��Ǹ�0.�_�l��@8����^���s�7;�����C� ڜ��A��E;<U/T���{*y��o�l��÷<U9Wzr�Ee\�O}U���]~���ݞ��,��zb�^��/A��C�]��N)��9=P輭��`�	
D�arA5�=r�H�����+�#�F�`�P�m�)��D2 eQ7l<�U��0<�XK�)u��t4c\Zh��i���UZ��.�/<�o͆�9{�ў,2�ᗿ��~�M���F9ڪ��K՜�Y�՝��UV��UK՝����Z���Z���Z���Z��Uj��U��Ugj����^���΍Yѫ:2�2�4Th��Q��uF��u�^�2��՜�Yջ}�7բ�EF��T����w��jї�v�[�j΍Yѫ>��ל��^s��}y������W���_����
�q>g���

�������FB#!���Dd"2c	;I�}����o���_}|M��7���_}|M�񓯌�|d��o���_	VY���������`D�#(Ĳ1_��FD���3����$����}����s�/��J����H�����Vp�TM��Q7p"n�������aG^Y~c�N��%&��v[�BIz֬�����kN����G���o�;˔�K�j]�M�� ���6�[_�^���x�[]�^��d�
G�Jp��[��衈T-��y#���������ܯ%�4�R���[��a�V���t�$(fK�bǁ(E�;��^*�W���n{*�F��{��3�o-�d�����cǭ�\u:�E�HQc����t��q҄��*�2U
d����������oK��.#����2�t�e��l�R�J@���-�1������-�x�t��[P5��g`-@��ޗMj#���[��c�������P��w���}��s���m�>�����7��½��ޜ���-\��}�+!�l��I2^d�ChPŶS�V"4�����d���!��H~���ހnx��}*ϥ��x���T���>�+���/\�pN-�Ф�\�ߖ���j��{�dvP�B�(�>M���SJ����i
Z�5+f[����YYj%J��/�Tr���=e����-����27�F�G1/��I�k����u=n����Pr�5Ga���15ܞR����;�k%��H�5����rڍf���HܮV'M��er�ݦҳ���9\�����b2���/���i��+����{���^�k�܇Z��1���eG/�Ƿ�:"��{��UG;�	UV���YC��e��X|�B�{'��r[���?��������PR�*P}E:����~Y�^��������[O��k2����|�d�vU�S+��j��S�*>�����:Գ��$\��"�����Ȥ���VҰ9yoKWr$�VU��^ʎG��*��e^���A��Tu{�~�GW�l���5�V�U�^�v@qM^�SW� ׀�ݐ{��j�qMX)��5}QM^�{w���G��0��;V�J�QIW�����zj;�*�/A��Tw>t~�K�Q��T�P�GJ��B�(^���t�z��/Q҅�:^���������z^��������(:P�O"��zj9��G�������^����.������N�ö�n���I��}R�����l�+64�o>��d+���,ܑ]�����r�s�S�-lk�����n��fµ.��͎�z�����y�cǛ�lw%�^su�Mj]���ۆ�l8f��_Fl9�f�W�9��Q����^���z�Î��V�_�����޾l2���WE�9���/9z��E:��N]}�J2�Xe�p���jիv�8g�^uh��;�}�h�v���Y�j��a�G���e�իv^��z7e���>��ל��^s��~nnnn���}ꂁA@��_`_`P^P^P^Q?�?�?ѐ��Dd"2��FB#!0�����$�>�a������_}�� �a;)�D�"V+)��Q���,��"��E�xXL�JE�F+�V*H�dJ�
vo��}�����O�"��B,��bY�eQ7Ⱦ�M�B,ௌ̓�J�n���Փ�Ұ�%����j��8���VS09z����B�(�lF���G8ڶM�Gk���Dj\T(?���vJ{^IO�����6���1�d�6���w���x�:~�+�!�M�����w$�WO�ݺ|��C2^!��m��qX���7O�aT,W�Z����P���~G�6�f'�#S��/�tB@�H�-��B��賊Cd)�2��dub���X�-�7X��:�4��V� �.A�.:B�.:B�.P�t��x�-�rPGJ��n))t��% Y�W������G��.MP�4X�d����Ϗ��<����)��fK�P�GI\�m"�Y��|b#�_mB���a���8>�,��Ӥ)�^! ?T[#��M�d3%�$s������Y4o�t⚽�6���B��z��Z;&�}��:�*���R�����<����[ Ql[�Jz|��D`9N������i�ܔ6?[��ܲ5l!0�%�՛
_��r�1����v�9R��5)K���.z��^��B���].4R��Ԥ|C������r��U?)��5��>l�~�:*[��!�K��--�x�\��S��ҭ�,��A�{d?������r�*V_�J�z#���i�������F��7�lF�c����:�F#{%I^ߗʕ��_\D� ��[8�l3]�K*��/Ӈe��c���r��&n�pli�=�=��G�jG��b͒�g끨.��;��NZ��\�r��os����*���z%�RY#�����<S���]��Ҳ$~˝@�XB�e�K$W��E|�$�}2M��$ܼ�"���4���%lvE�۬�yo��ʤ�VU%��>����ܨ�w*8:��Q��Tu{�_�W�l���3�Q�/T{K�Ҁ⚰SW���G��Q�/T{K���G��Q�/}����~�^����xa�/���l�A�)-�b�^*����ܨ���9�U�����^���t�z��/Q҅�:P�GJ��B�(^���t�z��/Q҅�:P�GK�S���e^�����W5<��*�j8ʍ������z�7/}�IP�Lm���+���{d�tw"�p�pzǮ�Gi�c�S,��y8�����C��n5��ǵ�vKz�6����Y�D��sƫE	�_VM��٪ߎ^�;Y��͚^��hյ/F��76��Do4oT��8�O79|y��V��g[J3a�F����Z��5�o?�󸻛D�枍th�k۳_69y㗞{�՝u�붕m1�cƵi�]/�/Vue��G��K��Q�w�}��:7Ωu|����R�gj�[��EV��n�/>��ל��^s��}y�������������Wޯ�_z��}ꂁA@��Q>g�q>g������3����|g��?�I��O���]���c	;��}����o��}�� �a;)�AN�%c��XA, �VVVRxD�'�I��M�ro���,�9<"Y�'���K!o��,�I���Dݯ�}'�'��a.ɣ*��Q�F_g��iF�c[�-�~^ߩ��S���8T�ƈG6��ʗdr�(�;80�~�"Z����v|\��R���k����8��B���P�۱�^|r��B�k�\n�j��iP�Z�/�W���j]���)�ީnJp��@I~I%�"�ㇿ��E��B@C=��@u./;~���~'^���{"�x��߮;z,W�⿐����U�B-�8ez�~-�aQl��HV $�CO�h��E�RqHl-�#����X��:�1J�X�+~6)e�K/��Y|l��g��H2�H\������P�Yġ�J�\Y��^�GYd) Ų:�ߑ������2���}7~G��W%ed���yB@~�/���q腲?S��\P;��*I����1���c�xoy�)��e~������Դ�?=8���A��L��D���/W�������K�8�/��pc��l��t��C�ӈ��\���./�T~5�v���(oܣ�}��4�Z&�u/|��ծ2u�'�[�2^|�(ԥ(�ą��~����퐣!0�u�ÿ��[��vd��Ί֛��i��iM��5�jΛ+��gk:��FC�R�:�JR��R��ѽ�l�؝�w'����=L���e=J֣�!���3Q�䈥�)l���[-6_c��������/��Vu�9#��ҫ9=:��ϟR����j^R��%m>��l����_vr��VScʧnnR�g}�1P;�|�.�/\Ų��j,Y%}?��йf�2,@C��<l��gż�����D��I�li�G|�<ՏKY����Y���k2z�������L���[Z�����,���7/J�trݜ���+���+g����v~��������!z�D/S���e^���C��P�>v����?�l���3�v����?�l���3�v����?�lυ�z������u�T���Y���d��C���<�[!����ew_�S���s�z��Q���9�>�����^���s�z|/A��T�^*���S�x�r�NU�ʼU9W����y�����v�)-]���p|Q[>�VEжk��l����{�����dx������������dS�����w�$1���V�U���!\��(�
��%I����z�6A�u�8a4�_m9�J�p�`u���E�B�
^��⫝̸��g57~�R��ݤiF;%���D�yƸ�y�����_V7C�3u�w�Z6��j��sƖK.>�Q͙k[�o��7j�[L8g/.�Vv���Y�=�yڻ�����Q��.ǎ�<,r�UR�UoQ�w�N�yu9u�L6��碌�]Q�v�yѫ:2��ל��^s��}y���������������Wޯ�_z��PP((O����O���3����|g��?��������'��?�I��K�0�����$�a'c	;I��X�X�X�X�,bV1���J6	��q�gc��7�<�,�}��~X0+?*��E����&x1�r,j��Kɾ�Q��FՑRU�DѰ�}��5�Wul�ʫ�ɾ��]��v�[�Z�s���W��\��nK%/rQ�J�t97N�_�`w���t��s�t*R��K�s��\�{�U#� ��Եe>D���`�)y>D��(��"7<��e����m�`]�f�N�d����۰�1���vJ�n.�o��8dq��99z�,��+�FGLҔa����߆9"�c�-�9!��$3����.R���o���_��ߑ�0�+��ȶK�E�_�@g0�%�~s@��_O��~�9��Yͷ��m�fV[b̎�ř�2��%e�ƕ��VS�iYM�8�cO�kn+X�d�c���{���S�a���)����%=�b9��Իd�\+�s�Т��m.?B��K_���#�������T>��Gr9��Ek��|L/]���0}��KL���Ճ��{v��tU��@y�-�|\���)&W�7H�0���z�_��𼏥���������ߖXqAZ�ާ`\GvU��&~�ݾE	F��e6��l��w9B#R��7;,�����'+���V�c���i/�g�ʔ��x)5�k-�ny�/�GE(5�>=%����A���*�J�Ԣ��/��T���� x��|p?���C�c���!�a�Xc�#�?%��=q�*V��]�E+�Z+�ݔ�WiPov���N�y��]�k�'�7�9R�R�|���>�M��}ڞ���l��Ȭy��žZ�S�P8��O�#i����%`��!������)�2%�ǃӮ|3\�t��K�"ϧ8��JT�,��c$��"�2���^�Ge�8�G�;a���8�K����H1���Ȟ^��֣%m>�������<��K$��&�e���&�m�oLVM�ɽ5��+g�����~ʞ/Q���80�G�A�{�2�}U�ʽ�W��*��e^���A�{�2�}U��A���nҮm�>*����"�[0=�̏MW����6�*�C���zP�W>����W�����{*9ʎG�����{*9ʎG������b�>���+����b�>����*�Hy��V�!�W2�����~��"��d�:��'��R��[σh;��g�=��;9z�G\���u��cc������1柷���٩��K^{-��z�����=�jŚ����$YL����=/��):�r��'nW��0����D�K<�9�j�iyK��Yt�.*:�*�!��uD�XhS�<�4�\�����'C�������o��%�W4�&~q�Ua��z�l�hھ�Yv,w]h�j�ˮ/u�>����~��Ue�m1�cµU����7W�N�.U%�q�枋O6��5Yz��^te�e�yϯ9��>��ל�󟛇����������ޯ�_z��_z��A@��PP(�3��8�3��8�3��8�3��8�3��8�3���6���|Γ�����}�%�O��RRRRRRB#>�>�>�>�!���Dg��|�c��g��o�����H���(�}�a	;I���&e���F0cg*���vE�}Y��6r�8'e�/�����v1����ܽ4��EЏH�1�g��_-[+�IdF)"����d�� ����<79?N�"��� 8v���X{*x�����C�޸|�Z��%�4�s�����?�s��|j�n{���r���s�1����JI��J�|	^�$��%z^���6寎/T>���w��	)$d@���W�rC;˔�����T-�䓵ܕ�����s���I;˔��ە዗����l�ߋd~���xd��?�@H��?�i�>����E��b�/��ȶK�E��+O�aZ|��tU�C��P:/�@~�l1����b)�����)�!�(<7����;^�K�S�����~-�V,��U����\�R�.E(�l��9N=�Џg�(ro��Q�~�g#FW()YY��e��jG{al��PvN^�|Z|�ދl�N�$��{��}��)�@"�\��F�H8�n�ū�,����n���[ӊ��2+�n�&�w�����򰽲�й�1�=7���|l��o)_,ss�Wc��e����VC�M�����ƨt���^V���;����Y����g=֥�A�y�q���^q��j6����b��������߯t���;��x�S�:G�t����Y��1܅�Ė���;�R�+��:�lddf�a����Q]�AFH�,G��B�-���� :�^+���4��:�x�ߊ��-Yʈg°$������|��2ӟ_rQ��[��#������+��:�����[�t�\/��R�;�o+�y���$�/��+>P2;����Ap>؟a��b`č�HН3�/$�����>
V��yx팭�XIjU}s!��O��培nY�������� ����zb�oNE�Ƚ�?eF��Q��Tl�z/A���8���B�^������FKOϕ��LVϹA�{�x>*|Q��#�0b�*��G�ߑ�ʡz�������"��dVU�ʽ�YW�+*�Ee^Ȭ���zm��~�߁��zm��~�߁��}���!����s!�J�o>����+�o|VO��=�ܞ��������%��0mF��l�trݜ]Յ⽞���[����:Zu@��C�62��{�~�q��W48��=�+5��E2����ǵ1���K�M�d����5�[m�3M
��H�[{/��T��+�m"�t����l���J�ʱ�iP�D����I�]�z�����U>V�I��,���@��ݠjᔿ!)ۙ����eR������� p���;S�.�E�
�Bϫ��-#3 �_�E���Za�f��ij]��^��+��G5UR�uTp��˿���.K��u���ל��^s��}y������W���_���PP(�3��?�_z��PP((O����O����O����O����O����O��u�gY�u�l�g�t���|o����o�o�o�o�o�o�d"2��������������ro�����?��97�ɣ1�"mW�U�����yI��<�<�`V}V}R��x�$����5�5=ll��ʺ;f�������P�<4.�'�A����e�e|�l��ǥ�z�aӏRt��8��='�ǰ=�̎�F��e�g�=��H�6���Z�Xpb���� �KP
��:E���`��#���Ee^�Z�`�!��N'�C�d���J΅R��[�%m���m����[׎C��K��]�O��G�VQ�iY ���K�-��Р��M�e�k�B�k�~��&ݒa��&ݕ�[��1r������'~�\0���p�?�I'��$��%8cnW�rw��}�6����a��������t��N��)���z^��Rۋv�)_k�d���){������C�;��ّ�W�.u���R��Q��h2oeN���Bb���:�,�r�\*��z$�P|�P�3��{�O-�l�s�yl�ϯ���C���r�E��@�p�n�;�*l���+�q#��/���t�����$�E�Tn�<ߵ�qz�R���T����Їӽp���J��e��l7�23���Y}��K��R�iFF���E2ߗ���DW������$P�E�[�E$:}���{w�M�w)���]ݎ'Q�;�Owc��bd9n;l�Ң�J.�J�Hu���+K�T�w�k�C�ķO�TiP�eO��Y�P�t8�Bz��&�������9-��`����¹͆k8+���/��������"P��ɬ�X�
�G�r�9�>�����P�߫�\�|ǒ�,����[)�2<i&�%��,LCN�-�R���f�{\on3��)�����̈́%@���?<~R��u��^H�+k_yz�d����h팭�XJ�u���W�jU}s-��2ݍs-��2ݏ��'�k��6�,�k��LVM�ɽ1Y7�+&�T�^*���S�x�r/NE�ȼU9�+���%P���+iR�6�����*6~��G-ү����x?���S��Tl�59��"�El�U�w�]��Wp|U�w�]����=6�M��o����=6�M��o��[�=2�-ʥl��+m��߃�ɽ�Y<Q�@u97����g��r�[J��m�}�U�vB�=^�Ow�A���u|1�.��o/o���YW�yݓE2��k����T��5<�/��㩙����F�r�6��@;�j�� ���{"��(�ơ�h��GT��E�nN�i(zhL�'"��Z�!���>�VFՇ���ͤ�k����~>�N��dZ�����g�BL�뷵�o��Q����9�F�R��*��Ȍm�hȖs�qF�i������'H:���Hn~=�6۴��z��.31�s�͍�
_
^]/.��wp���%�I|*7��玍�7��p����>��ל��^s��~nn�3���$���'��|�3�������
��D��O����O����O����O����O����M�&��q�g�q�7���|o����o����o����o�o�g���n�����������g���_g"�9g���(�BU���I	VYjO�Y/&��U~�k�ſ^�B�Q
E�m�%,�ӆ�^ێ�%h�l|�5|��{ ��RY�`�V�|�j=	С��Pa:t��I܊��봝�'z���|�1>�lS����7/o����=*Yܶ`w(rϝ'�������dg��жFpc�<��_Ǥ�mv���X�b�o�FM��I�1KR&� ��C�#��/O�b�|���㣻�Z����w�4(vr)*�ǥPS��KW;>�?>-�׎C�%�s�U�`�`�%/"��ϡms�[\�Ok�)�ue=�d��ݒv��N�rS�\��k�Gk�B��Y){�*��
��B��|vJ�-��e㲅sܲC�l��؍�v#��Եez���R��|`t ����A���V�ɤ���Q��a �ts#@�r4)Y��z!7��� ��G���3�_�p>>֗��x�g����G��KQbS�C1Ο����mv�Y+ٯ����J���k�����Wr]
^ˣ��%m�ö:��F���ѓ�����|S|Q���ރ��8;�Q�:8����В�j��`��q{��C�C�$�%���e>H�W}
g�/O�I[t����Z�f�n�G�1_��vJ�Ti�J�z��ԫ�|;yn��rx��RF��4���V�]�f�-���Zܶ#��e7�g+-��I]�N�)n�[���������D���b�����T������9���:+�����_�"���>�e7c���b��*A��y&Z��M�T)�||��Yēd��y-�|wK������x`˃����4?{�o��l���=}��_��8�u��`������$n~3GG��+d�-Z�\֡?u�)-Z����^;c��ly{u�/J���8�--��in6��`�����2ܟ�-��V�g��,�[����]�{+�oevM�ɽ��7��&�k�H��i��*�m�0�V�����eRZ����y���%���6�*�Tl�U9dS����V����El�Q[?V����El�Q[?MvE�Ƚ5���"��d^���]�zk�/NE�ȿq\^+*�ⲩ-����P�NY������C��ǻ=�=/�*��o����`8��-ʼV���wK�-��Ⲯ�O"���1]/T;��S�tq�_Ww�A���ePSW���Pw%���&�14�Z�r��;�}��핵�RHȮ�\��)ˏ�5yx�6�J�h�)����!d�&�@.^*gG-��j�˥�k�۔��P::��]�p4�+���{�<���ڊ�!6�)f+Y��W/���خ���f��l��6�si)q�W���+�?*lb���*2����vz�,M^���'�W�,a�/7|��N^��e陼r��� `n�Ƹ̉����Yrk��hڻF��{W�ڿ�9��>��ל��^s�p�p����o����o��|g��a.��]����
��D��O����

��A@��PP((M�&�p��8γ��8��`o��8�3��8�3��8�3����}'��|�_�_�,��B%��E�A%�g_���l>Ѱ�|�g��ݓ���h�\Xu��~T[
MY����0췜W/"��/�W�C��jr�V������}U�����tw+��{?|W���I�W�hu�:�z���S�����~���O�n��#��?�q�Ҭ;��8^�cܩ�z�R�z'�C�ި����(��8�or�I%��>�]��Tk�6�H�z
#��@�!��|l����;͔�Ge�|0z������R�%�ez�,��ro}Y܊Rw��L;-���QI7z,�ä���Q��KU)dr�"�jR(��9��԰b0yU���d��ЪZ�J��F�(��b0}�%K^#���Y!�H~E��d��DaҨ�:U�`� 1Ȥ�9 ���$Ҍ�Q���?΄��]��e�eO�l���e�*3��Fx��Q�9��CV����Qc�@K ]�:�{��7���;�+k�2�E$�������_����?{�d����w�s�7uy4�eQ��W/*e6Y���>6����p�,]��jv�R�M�8l"yߎ�����_��X��;`8=c�R�{�K-s]�w ���'�qv�:7{%Y��-�+��E2U��/���L��nyJ�w[ݑ����j;C�����%�Tʞ_�O�ۣ��.�o�P�p�|;y���K~OaO�H�ܑY��}Gwi#gr������d��-6'c��|�4�O��$l-�7�F�v���t;d;__l�������l��ƣSԣ���}?;m��GڰU}�I���u��YO�㢵�]f�ቷm)��'�V=�R@J=��|hj����s������|Pn��)^܁I0̭�g6�\W-a�BT�}w��r;�q�{`|o�1���+: �S7�L���9�jds$y�֡?u�*����::}'G���Ԝ��+e��[!�~�:O�*���������2ܟ�-��2ܟ�o�x����Y��<V�g��,�[埻}��OȨ�)-!�ze�^�����6�[o�r��*�+��r<U<eFM�����}so��b�oMvE�Ƚ5���"��d^���]�x��~(���+g�����~(���+g�ȼU9g��,��;>>+*���VU�����r/|VO����·���{+��Ȯ���ܠ�W4�^+�ӡ�t�:�:�r+"�Tp>v��ݾ��Q׀�~+~Gr��ЊJ��Y?�=��S#{�Yr+"���>q�.�[���<��L��b�8�-�b��:;�%�;}-?"Vbe����M���xJOeG#�����KEe^<�_��pd�GrKE{%mw_�Q��뻐���*��3K��2>u(���!���u�H��@"�[��ۤ��b��%�H�m�}���/��;Yڮ�9���v�t*�����%�Rf}#J��b��F@�:�41�K�Z����'�W�`ƮR�R.�07WS����y�34fu�>��ל��^s��~nn���ꄁ�

�q>g�p]g�p]g�p]g�p]g�p]g�p]g�p]g�p]gp��D�#:�3��:�6���W+�OTOTOTd
3�'���M94L�J�E|"O��'����Dl�Q7�İbZQ��ƿ��J/���0�u1�����dp5��YO���7�r��	[J�������!{�^���]�܊��En=U>~��oUO7r�����T�=�^�����W��+�o�Ш���7�~h6���|���f��V<|�+e��mv������:�>������ǿ�vϰm�ρZ��G_M��-�t�1��$̵l����|�p��q���gcx��禇r��d��YF��S���?8�|/Q��ǣ:ȌzOB�I�
�\:�Z�W����:�������u�������t����!�)j"���%t����ó�vG�-C���9F&�ä�t�#��1K]7�S���b}v��j�,�푾��'�+��S��P�=U8H6���q�����Hr*�_C��Et��[��x�-��ر�Ŋ��x<|,�|>�[ ^43�UP����h����Rԏ�C���K?��[xs�-}����� �I"��e}��
���8���C���;|����IX��8��a�������+�G����+�c�l���oo�K}ݦm�l{��{e.��Ee��dd���6{�M�=��l#��+g��Tj;[eGy���vs�~�Y#�|�k��-�z��T�_�VTm��}j� ��v��VA�C�{̾�;��m,��fV���H^������r�ϕkS������FF�-�0��.K�}����|����S=�ʌw-[�6����12�+
�ۥU�W�����e+��C}��f�ۯ��G��ZX�J|�d�-i�|[� ,�)FZ�G:~�O���J��rKr�e���^��A�J�������v�����XH�E'���9���|}gGY���B{)T��>7���tu��;c�۩::TL���k�&��F�6��*��J��Ҭ ��������]�{+�oevM�ɽ��7��&�Wd�mwGs��!����^����W2�J���Z+*��p}59��,�T�*���S�x�r/NE�ȼU9��"�T�^*���S�{*6~ʍ���g���*6~ʍ���g���"�<|�%�ae*E������1n�@pUU�ʽT<��K�Q��Tu�U_UGW�A��P{>u�UO_�Q���t�t�g�ʽT<��G?�S������UEܠȽ�eG�A�xj2.�G�Q���t�1](6�&��>��D���::Wes]�{�{�+~��`J���+�+iXv������nY%�9<]��k���*���T����l��\�y�[��뻜�wrKE{?q]LWK�Qȅ�y�O"��Ik~�/]���~N!(6�>_�S����s���)���i�NU��dPl;KǮ�H���j���>7�M�s�m�ү���p�̌��oi��RV�^N߂�UW4�?��;�t&e|��^s��}yϯ9��?77�_���B@�
��8�3��8.���8.���8.���8.���8.���8.���8.���8.���D�"n�g�q�g|l�W+�OTOTd
2����B+�ѾQ��x��T�udV�e�{+ڴ���zې�7
�m�폩�=���rt�<vO��u�*3��D�jT�[�����������%�����C����-�;���w4/]��v��n�-����~���r�?ܷ���x�T}Q\>��s!ѕ�:��V�q_m^>����l�q\�q�k�}�����߆���}�Σq��������e3A��Od�q�tKT>rղ�C�����~��U���I��I?Y҃k��*�or�σ�����>��$/Q���?�b�e�dF�I-E)=p�\3� ���#=p�\'� ���"x0��:7� ������Z�W�QIg���`z�/\Y-@+�0F(ã81H)F��G!��'�C�����^����B��W4�~�G����㰞Ȭ����G�d��Z�#����f)zpm��<7��o�������+�0��A����G~I�r��G���n�%!b(�6�(mܸl~��k�5;��=��m�E$TR�ܡ�!z�oN=�Р��-�]?_����q�6�f��~�;��o�O��%�g�S�=+-��P�[=���2�*�����I�$X��$iݵ����FC���r>��P�xOk\R�:G��Y�� �tzC�T�=�ݼ���6�dw-�d�vH�ֶ�J���v�*1C�g=��-�yn���5�k�l�������)*��%���'�����
�i++�I[K��1�y�i@��e�*�������	>K}���o���~U�fƷ�J��jT������=�_�ҳ�x��g�VVm}�o���=�d���������^VԶu������I�đIl��d�����q�=gD��s�k]`�|%sZ��i�>���Xq��N��I�Ңk�&���r'�a��X~�Vl�_�u�l�_������]�{+�oevM�ɽ��7��&���8����iA�ܫ�]���e^�~s!����9-]Ȓ�\LV��S�B�</S�B�Y��"�Tl��?eF��Q��Tl��?eF��Q���8���B�^���p!z/A��Td�*���I�fN����d�nV�u}�^�#�l�w(y�����ܠ�z�:^��΃���|�;������@t�g�`xhr�U#�Q���s���EܠȽ�e�A�xh2n�G�Q������<�#���[5���/���w}U�/|�����5�X6����{�z^������x>����+g����벯ݿ#�o����$��JKEu�OK���T��z�Gr�����*8=��/Q���wz;~�]�x?�v�Y)k�<�|����7��Wu`���Y���>P{;�[}��"fҁk)����}���6ї��6�LL�a%���<G�/�ג�)K'��XuU�Å�_p�_N��ל��^s��}yϯ9��y�y������
��D��ۇۇۇۇۇۇۇۄY�u�Y�u�Y�u�Y�u�M�&��q�g��8�3��8�����d
2��I�_�Y��'��a��'�5�We��p#ZU����m�4�G;F��ǊIed��G�p���:�O����Z�ֹ��d;U̇k�!���xr܇��!��ҭ{-�=��~��?e�G�ݣ�n�\ұ�4�|�v�/n�+c�em����:攮iH6��۞��ܽ)��n�6�>=2^K�bݢR�q��-o�sox�����^C�������m�}6��4�a�k2�F��}|R?|�V���j8�����Hq;�m'�"�v~<��+m��v�A����徾�n�-�{"�}��U�z��Q�Р�t(�?�
���B��l�жy�[<�����d'z���l���#=v��������ǩ:q�ބz����<�b�x0p��8^[�/]�����;e�r���o�$g�#%m>_�]���x5��6ӝ�B�Q�D���|���oN�rƟ(����h]9F�����s���}��G�����P3d���>�_��g)����$�T)�۹[ݕj��_z��<�DC�s��`~�G��Q���8}�=΅�o�S��Puz:�G�Q��7(ˊ�&�>�$/l����^)�����C�[6u��_��⪞�ӡ�yY��ޟ�+ag�*�K#�g����m���X��=>��I<��$��?�T?��Qf� $����R�/��0����@�������|�;��7�:�g=/K%�g�#���3�>s#��;��9~�����Z�g�j0����s+?!Q|����^&ͷo�[��1Z�3�C��6��싊�o�����_�|�������o�B�V��A�⵪v�ۯ��rP�:��2��WzY5��m�)�z>^������u�Է����zF�����=�/rG��z�t�Wy���2�k��\W/�d�`�2��<�����|������t�N��a��ly{u'/n��d8�6C���t�l�c�v0l�c��zm��}���_������*���_������*�|o�tr/!�x��|VU��w+�0l��+d;86+��p=�?}Y��=�7��g����v~����Q�{�2o}FM�ɽ�7��&����t;?���C�����t;?���C��m�n���/]܆7����ϗ���m�5�W?�l��G�;���{#���ǲ ;fDl��[5�t���Q��T��U_U#�A��[0=T9W����ʾtW΃�ܡɡz��A��Tp{�97��&��8ʎG������7=�K�#�t�:����λ������?}OvV�y򶕁���(z^ʎ�+g���*8>ʎ������b�^����+�����5>�棫����/}G?�Q���s�u�}G?�C݅�.>[�g�S�r��v�V��VH|>��C���u}T.�r�o�w8l?e�����H�؈6'"GK}�uFn�RH[��;^��f���JWr���u����<~����X<�RyI�9#[(m�w[�ל��^s��}yϯ9��y�y�y������
��}�}�}�}�}�}�}�}�Au�Y�u�Y�u�Y�u�Y��#:�3�� Q�g�q�gI���d
7�7ʓ������������#q�X����&��,�YĤ_[�lG)("�;��f_��a���rZ+�V�xx�u^�|��]���u��
攮iJ攮iJ��9[J���NV�h���Pl���1�2F9[Z����q��\|v^V�����:�򶞮c�6:�c�6���U͹+mΎ��kOH����#�/�W����iN�Cr����?q��?�u+i�-�sJ����B̝^QVH�d��4n��O�n��C���������O�RA�l�XJ�͟�L�������}v��J���s�Ү?r?M�7�����ܮ��Ws|�>q]8���WG�+�������q��y�U>~��8��������j~|5?0�A�����y�t��N���C�(���cֽ�;�l�86C�%�Wz:��c(����2މ-n��p�d$VP�Vw���S�v�O��)'��]O�����������1c��������8����g�����;�n�J]��h���f��Gʱ,�-��^�@���?res$W��E��[����<Rޗ����d]
����H��:����^���u�r�el�
��+���bi����1Z�K�r��2��ϳ#?)�S=�D�C�FBa�+e������w-A���j;���#�:v;o�Ej0
�z�!�m�w��Eh0��%��h<z)R��)q�w=�Wj6�H���QI�A�Kr�N�Z�H���>=n��i��kL.���Kv��^�q��؛����햱��b�|�Z���+�-����ʷ\�p�[Z��k�����\��yyoGbd]9/��Su�l|ۻ�>U�B��D?pb���<2?k���m��J|����|V+ơǡ����vC�o�烊��d��Hv��2C�N������t��	[J���G�-��ֺ�)Q?�tg/n���<��O+m��*7�!��d8�e���o����=6�v��]��Ed�Ȭ����"�dVO����Y?�+'�Ed����V�vuͿ�S��Tp<5�W�o��e�������(2/UM�ɽT���ܨ���8?:�·g����v:�·g���q�=�ǰ`8�����0{�d{�x�K��������O-�(^����;��^�{#���E0{�L�{���ǰ|1���^��|�=�G��Q��P�;��T����>���C���e^���"��/M�A��P������{*9�����-C�,��~�N����z�{�:�rC��Et�QK� ����䵾��ʽ�6�"��2�^�*��2�^����x�z�mO���W5X6���t�U(^����{�z^������ܶnw"��}�W���J�%K[�"G�T=�L��P<P�^��ܨ��+�]��r��G��v������d����8k�+�����*�H8�Qyyoc,�ԮI[A��G�z�N�S,n|�� �O�[��n�P��~�
��u�>��ל��^s��~nnnnnnz��A@��_nnnnnnnn]g�p]g�p]g�p]g�q�(�d
7��|Γ������������c�c�a:��� n��*�/*��*��|cr��"b;[-�=��q#c��Ux�m��n�ܕ��/Or��/r��/x2C��+�rVے�:��Ύ:��>������J�~R_��K�9I�W��U�)�|	"�$_�֧����I-O~��M=駤�u��Ҷ:���8Y#!ef�F��I���x6�r��/$O��'+i�^�����Z����c���af�׃L���k��6����GZ�#��~&�ʁ��+RW�Y�����(6�q�\zc���N_�����䵺_�J��Q�Hw`��!��Hu}�_|�W�!���u}��|�G�-��[��%�~�/����9o7�ߣ�o����Wmw"�}U:�8�ߜV�Χr+?��r�F���[��r�-n��ְ�Iݺ8���gn��PR:;m�g2��t�
S��宄�aeJK�á���:\���=qf��JJq�b@JqlX���-�q���&P��ȁ�X�ϠY��D��H��ܙ�5~=v?�G�U�)-O��֫�R݇��'��5sn�W6�W�����v���I��v�[ׄ�{4�\�j[>/ݾ�%�1c)(g5�G#�����oEq�����͚^�&?���sf��F�U(��_n4h���2

&
ϟ�a# ��`�i>�}��I	���$lp8mBs����G;��n-a�j�<2�j��/�^^⬿[�D��k�6���%�{
��x��0�,	ec^U�I�/)H1ݞ��l8�ҁq��--�$�?>��~�_ew#�oȮe���;%L�~W�_�+[��w���+c���ߝs镽/K���W��� %~[��4/B,�2M���<z�+d��Q��C�:X�Go�b{){	V+���i�oH������|������Td���$�*�Vҥ�̇'�d:�^C���H^�_�k�z��+'��d�����S�w*r�|VO����Y?�+'��d�������+�oݾM����2n�ϡA���v}��-���T/C���$P�MӡȺt>�FU�e^���l��[0=V�U��l��[0=V�=�ǰ`8�����0{�`�q�j��q|�7(Y��g?)�#j��|�8��r٫�dw"�=Ȧ�=��`���=�f�=*�ǳ��w�A��P���/}�U�`���?8�Gr�*�[%]�f��"��/���t9l�|�80�?�Q҅�9�����G�~u�dWK�A����~q\�^-�l�g8��8u�K[���N΅�r�ʻ��Wr�*�[%^�G������j;����A҃h:PmK�Q��Tt�z��/SՅ�z��~D/A��E9+��d���{!��:F���11s#W� 0mr��xm�~��g�C��Ҵ�;g'���܏o�	[Q�h{�Z��\�u|;Xo������bF��h;����\�1M�j��Xx��><�_+)�;�#>VT�YL	YZ�~��1e��}yϯ9��>��ל��<� y�y��<�!.z��}����������8.���8.���8.���8.���F@�|�7��?�?�?�?�a'c	;�)�AN�
u�7��o�FZ�}�����j�D$L���C��;̿9$f�m�|	�ҝ)�ۜ}i�֜�=��Ҷ:��ԭ��m��֝i�֞i$��HA�d�č81Y�+7|	�#O����eQ)��i����䄭�+�!\�
�Hr���<!��������q7�2E�F��Lx��ZA�!2�1#NH������Uyz�81������̾i[$@�25�>�sOx23��Z�2�`�zm�.�)D�y7��u�V��zԿ/Y��l%�Y#7�Z������Lu���zS�� �t�Q��Q��V�����[��O�n�������v�Q����_�J��a��u}��}��}��^[B���!���b\|�����z�_)/��*�*2��kk�����$�3���[�M$�*���9-�����-���s�B��=�Ǯ|Y+{��_�-D|?�O��5͖�~��&�R����k�E���Z�Z){����gP2v�f��Z���v�NOީ��m��}2ã��zm��U��&�+5��?[ׄ�uj���I|���C��8�(1 ���+S����)m%ڲ��X�BUQ���D�с'��qo�qoܹ-��ī#_WV����i��b�(S�غ�7��;h�:?�B��5�;3�Yy��,�9d�Oc��Ŭwg9yߣ8�4K�»Uw�dĲƓ		/FǮn�e�����&�������/�9���M����d�w������~����E(-�?J�V3�~�2$Ron�g��r�v��q��~?�s��|v)����{��$E��똶Z����s��$w��D}<,HG8�m�����/,�2q�Z;I��|Ɒ�������ܷ,�e���&���ϝvO����|VO����9gr�,��d�:���Q�|�2o�FM�ɾu7Σ&��d�:���Q�A�9?��,�Pd��e��gӨȻ��?evEܶJ����ϡ�w��}�z��Р�t�{�`�q�=�ǰ`8����%^����xb��RU�J�1IWB)�d����l��dV�P)�������cܞ�f��)��g������=��g�m���U-@%^�f�������(z��f�r=��g�"�?8�G�=�ܶJ���|z��H�z��gӶI�v�7·g�ʡz|/A�{�x�"��p}�<LWK�l���5}T9W����z�Y�$/�w��K=�̈��ȽV�U��l��[%^��������h:����ّ��{(:���������*;��~��+�ܶn{�{�+f��r���6�+�������^���rٹއ�����Ȯ�l���.]ʎ�������hz���/݀��^����)�Թ �~�GC���7}_=�'��ܩ�~�9������6�l;��R��M�}K�յ�u�>��ל��^s��~nn<�<�<�n��_z��BsBs�'9�s�'9�s�'9�s�[�]n�u���[�]n�u��q�g���I�I�c�c�a;)�AN�
u񓯌��6�de��t�/�I�K���-�ڵ������S*�����:�Zx��Q��9~��|�Q�$���?(�)�>H�/�� �Q2�1�xG��t�G��x3���������$g�#<	�H�Fx23�����������č8Y�T
���U�2wxB{n��F�1Y�$i��bS1�H��18|��@��	��%��4,�f�6xx�i[L�13�������$gY͊�`�<�Wn�Ub2H�K1\�'Gn��N��<��I!ej�GOA�׊������[��:�i�6��i�6��c�6:�c�M��=1׊�?v�v�dv��;W�n��_�=��/nB�犔��^�u�^C��h�rv�M������Vj$���BȥB��څ���y~��!g���b>���x�����"S�ao��d��8>�����X��'%giڽ��^̗�n"?��ȉ�V��
���ߕ����%x�6/#Rt�x?�e���Iܧ�z��Pw�/O��kT�jY+X̷��Xw-��1Y���l�����n'{b�� ���ql���7srYI��v��Y�2iuX���E��dލ�O�\A�o��)�.��c�O-��oIB�ӴY���ڂ�a�2��
����eB�T.B@B�ȏ�V����
�VJ�1\Cs+*)#�
�G���6s ��#����[���u~�;��իW�"U��[�oH���D7�-��o{��ovuLw����~���*������T�Aᖪ;}:+�C�GvU��E�\��,i �;�wi��5�#a���v8���a��I��:[�㸝�g����6:��+۬�S;�����I�D�'��l$~�[�^*���Q��T�>u:O}N����k�/LW���+�~����&�Ee�ʜ��S�|�2o�FM�ɽT��"�Pd^���A�z�2/UE�ȽTr�"�Td����l�w��.ϡA����V����ǰzqK>�R�����0}t^�W��x`>���`�`>���0 8����S�`@qL�R�#s�t�4��N�\��k�os�C����}Q�/TS?���G��6���A���4���Z�it-���gr���5ax�G�)��J�q쏜{#���G���I�)"�[0=V���EޏK<6�>�U��{�y�NY��]�f����t�x�d��ǰ~t=_TS����9�mw�Ƚ1Y4]��[0<6�?���l��P�=�=/eG_�A���%^����*���=�_}W�Q���u��M�#�C׀���U�g���̷_���!�^��獵��n@p�(^=�܀iw�[���N��d{�2�;s���ù 8s�r��7r���ܮhy��K����8|T=�^����{#ݟ?��}�#���x�}�}G"KP�}���^w��>��ל��^s��~n<�<�<�n�З��.h-��8-��8Ns��8Ns��v��.�`�݂�v��.�`��7�7�7��I��X�X�+���I4L�ы8�jUȤjƢ�W}��e�:���mǏ$@��o��#9y"|�v}v�$_��'��.�9J�<��ǦK��J�%#�	Y�p8�KYA�pc(�4�	}.R}.R}.R~�>���k*�YT
ʠV],���ɺ\Jb\vM1/P�5�P��������O��]�6;/FGl���G��P15jf�FT��VP�'vj-B�L�q�qؔ�c�vk���/ek����z]C�����zY���#�m҆�CUO�dT}r^����ђؗ�t�ڰ�/�S1��}ގ:�֞�!%��@��u�֒ZHIi!%����Z���BKV�mi\֐mi���Z��]�S����}�ڰ�v�^;|/��:��^�깧�m1+d�<|�k��c�=�����B��H��Bޝ@�A��������}>���)��f@z��%P�����_��������zW�څ�I~R���V2hT�P����!]��9?�y��͢��v��[�*6_C��Kv};}�/#u�Kt�;td/Z��!>t���t�;+i���>M���}6�g�C���r/�m������7d�2ݒ��|�����+a�v�
�ǇY!H\�˓���5��$]UTy���'+-���:V��S���ŞY�N��@����A��7����dA��e ��Y�M,���D@Eӏ��t�?,���M N<���zs�Pj-�����r��hR�H��x2�Db���)�z}��[�d�����N��G�8���3�^�78(�Fa���&�?�'��Fjb���K�N��#>�[�j4�-J���k��9l��h}�}7��ʧ�)�kz4BhHN{T�-֫;FJ�B�����<�o�5��T��kE|�9v�m+2���}�l��Ҡ����\Y����9g�+g�ʽ�YW���ө�t�2/TVYܩ�>u7Σ&�Pd^���A�z�2(�g���:�C���vp����t9��'�P���MފY���}:��Q�B�Y�)*��0z\E��`pb�>���=�ЊJ�0�S����0=p������?8�G�=��d@v̈=�ӏ`w��n�R��F�W=.��r�������~��g�it#�����=���xh;�����d�`� =覗����v|흝�f�r=��g����{�`�qLTzE܊H��Irف�Y�����zY�Y�-��d��l�|�/� ��P�}6̈^������	F�����>����Ԯ]�d���@q�U��l���0=V�UUܠ�{�:���r�*�[0;���U��{�z^������n���}G?� ��Tl��7B�އ�t⚼}��lׅ�9�ȧg�ّ�l�p��Y���0��RU���b��;gdȃjr�U��~�r/S"�q{ ��w#���뻞(�l/����*O�J��;���"��j��[z1�Ff��z'�D�9�ם�yϞg<ˍ�7<�	�������p��BsBsBs}�ꄁ�$�Q�ѿV*���F�c;��M�Xϲ���O}���H�G��"�e|ln⸜ҳ'�8���5�~��VH�Y#!d���3���uf�:�#_�Vg�Vg�Vg�Vg�Vg�Vg������c81�TL�|������\��|��L�ɡf%1.�2n�P�u�vef^��QvK�U.��Y�p8�s�g;�v��)�Êj0��<�_��]�2��]%�iY�xʽ-2^Gl.��EYY�#K��<�o�FS2٤wGL�P)��>M���d��9=�b�MV��테?/�K�.<W9[Y����h��8`�j��#:Zˣ�+�e1#Ne<��G#O��������i��3�����Ώ&�k.^�>^�9[#_+dk�l�|����dk���):�(��C��9z�V�^e��㽳�r~6t�]f��S��G�pl����_B@z�6N竹����K ځ�����W���J2�+�2^Gb�ռ�<��K^J�V�1�d��G�MU�}�y{�b���&�E䴇I���i�)#Οk�Z�%��z<��-L��V����V�Oܑ��n�zd<�ܷr�~Yt�!b9"a/a����A�B�t�Ѓg-(BM����e��,�w�R�$lf��f3��
ĵ��H�d���0`ϧh���c4��	�%囖~�H�:�(	�"4�n@�N�p�D@C ~D��� ���:�283uI���:嚡��3��:-��%P�
8�� VI'��(U�ܡKQ�Pug�A���$��|^���%�Q��5��8n&���ͫp�AQ�[y+�Eڵj����g}��G��N��0�)带[�Q����~ύ���e��FڻV^�8p������+Q���������$��P0�mc�;�j՗���n*��ڈ�X1]�x�<?�t����IgB�cӠ�=T7r���p}�W΃*�P�]
N�"���]:��C�t�r.�EӡȺt9B�gжY�-�}e�B�gжY�-�~e���,�Ԩ�)��H�1�z����`0S�Y�p	7N&��$�8��N)gӏ`x`=���(�0#��4r=&���n����]�t��/TS��Q��C�%}�����$]Ȥ�� �z���Gr����{�z]�GB����z������=��k��=�
���KW=^�{vKT��Q��|{_�S��Tp%���S���l�t���t"�|zM��!z��C�w(r��Yܡ�!z��ȡz����G����/l���x>�/A�B�r��ܨ�w*8��Q��Tp;��G�Q��Tp;���A�|�2��K�C��[%]�frفܶ`w-���UܶJ���W�������x>���g����v~����*��e^���A�B�T/A�B�T/C���8���B�^���paz�G������z�/lՅ횾+f��٫�j���z惥�����:���l��[5|V�_d{^����4<�懟\���c��sљ�D���;��;��s̸и���~y��9�s}�������p���ꌁF@��Q>g�q?�k2��F,`�0I<L�ԓȱ��`ձqR6�
��!�ߣY�]��3��Ǒ���ʼNx�]�bP�)G����Vo�7�՛����uf�:�#_#�l�&��4�ɤvM#�n�����x�,ĸKɸJb\v%%�)/�x��}��;P�ڄ,�_P=�xE\W�W�����O��<���%f�%��/9/��%�q\������yY��be�|M.��7dv^�/�b��5/C����y�u0���g�e��h��7�3k�C��7��ц�Pe)ǳ���޵,��Y͜d��M�� �v��h1L�Yx�7�Ytu��b�G�ɡd����������d��2w�;���N�1�������������7yz��^�vV��d�N���ݒ�;��)>����Or���x22j'�֬c��]x��]�	5w^۷�)E�)BP��\�JR��r��f�g���r�o��e��r��6?�r���Yhye��m�%�l�WXfL��?�p�v&�p�k�}�;��;��1��{��R�����Ar��(6���n�����zT��-�W6������򖧆6
�4��Q�S��?r:G�v��4n��̬��8�&a�7�r��?i9%R-�N�4e$n�M�����w�HӉ�7I����e��cN�:K�X	s-C83��:�N�	2��垡�����ӆF�0f $�˧�9�N�YtထkN�8����1�RiçRi�B�j
Q�@_z@Ih7�����
�i��^�{=RL������YO�ָ�Z_q�m�Ev�\�ʑ��f�[ױ�vJ�:����GҶ^�ˡ �z�տMG~@~�+%�A��J^(>Ο�pl�%��F�V��ͣi5|omˋ	΍XK�=|�U͏<�mK�u������l���T����z�����`С�|���'���_:��*�P�=T9WB�*�P�:t9N�"���]:��C�t�r.�EӡȺ�>��ϡl��[,��>��ϡl��[,�T4��D�qLTz��`t��>��$���pR��Y�p	4 �@p	4 �@qK?� ���0e��=&�E%����l��El�q�/LWo�!��h|����"�P��������[0<49W���ܡ�{�y�d��Q��P�=v��RU�g�-����N�����Z棫�Kym�����p:u<]V��t�2.SZ�W��>����A�B�94/l�B��d/l�B��d/C�B�94/C�{�/}�E�H�z��Ƚ�7��&�Td�����Q�{�2o}FM����v~�����g����x��r��ܨ���2��U����x>���������x>���������^�"��8�E�p!z���B�}�A�{�2�}U�ʽ�W��*��eP�G����^���paz�/Q���8>ʞ������j9��G���~�8?��EsCϮhy��?�C����tx6ٯ�s��|A���r4fh�љ�D�4O�;��^s�иЁЁ��p�p�����9��>��_z� Q�V0+��*����<"O	;�	y������Wɠ�����G����#���,���a[Kz�p��)���֭t��\�G9�1_�GjvR�)��)��)��)��)��)��)��)����%f�#�	�H�BGjơ���ǵ�{Y��%��`��,�8jG��?`�~N;��q�TBwg�wn�?+�om�6]�l�]#�֡%�	�I}�����U�z0����vԗ���?)~��be�g��Ck�@7���چ2֫U�.�q����Yx���\jճev=��l�]���F��
+�����\bsH���~��m�aL��VX�%�eг.���z=E_P���@�ΠbgP13���L�&pc81����x���bg��g�����w�y;��E�N��'GYq�GLq��G$+�{���}�V��<��^o�Z(��Iyߚ^��7j�Mg��>�o��_sM!P;i���X��Hr�o_{�f&]��������~z��0m��S��kW�#�Ο����G�^�\�`��/��[�}���^C���r=�=����eO��v9{�1ڮ"�?k䰄��F[��>���܆$>5gM�e�RV.^^^Oac��z]���H��:r��DF��Ž�@M�Dp���7��X='r��|��C-;� i��'@EӍ z�i�*H�1�<��;�"$A����4��5�AӉ�\����h3:w�Knpf�"�MoN,A��~@T��c������9&@�o-ӴY��s��Y+�7���e�l2=���K^�o�V��Կ����=K�e���R�*H���8+R^���C��8~"9gax�^#� �4�JZ�e|U-mk� �I�0ݵF�l8�a�_G2�$�<M%��Mn���Q�ͣ��E�4��N��Kể_�k$V���\�xazg)�B��Y!��]7��t-�~��C��P�<49Wz�*��0z�>��ϡl��[,��>��ϡl��[,��>��ϡl��[,��>��ϡl��[,�TJ��E%^fN=�ހJ�R�'N=�ӏ`t��8�N)gӊY��}8����@0}P�{���G�ҍ�Y޶H�6�?eG�ntt��1$d{�{��f�N�"��d�8��=�޶dw��:�ٟ܏d|��:���C�w��~e�rفܶ`@tO���v���C��R�G?����p:u<�*��r 8�S�t�u�e���,�P�����A�{�2�}Y��=�7��&��d����Q�{�2o}N��ȡx���ȡz����!z�����z����!z����!z����!x���ȡx���S������;>�G�Q��Tl��<eF��S��Tl��<eF��S��Tl��<eF��S��Tl��<eF��Q��Tl��?eF��Q��Tl��?eF��Q��Tl��?eF��Q��Tl��?eO������߃\�p+��s�W1Y��ɫ��sQ��j8����W4*惥�s�T9W�������љ�3���h�^w��>��q�q�����?������}o����(/(���D��M�&��A$PI���_&��Y�F0cn���դ��Iwn6{�mzP�kD�|W-|[wk��\H�efN�Y��dv+�b�$��8�Y�H�BGj;P�ڄ��$v�#��.�r�Y�b�v)�b�v)��)�b����?_'���}	�q���~�w�#���z�}	�B��k\v�#��w���3�C9�=�׻ڒ����^��{8>��Kg�������5�d�*�q�Üwj��-�u��_٠.p��_��m��~w��ȇ��̍����i�����%+�4���Xx���nJ� ���{s{���x��}����#���b���x�<~���{P�.��t,ˡf]2�Y�T��e�.�w��x���q���������9y�������x5��#<���ܐ��.��)��ڛ�ĝg�櫞:4jݣV�Yz4jݻ5���p��5c�R��dX��6�Όɗ��͆���Wߴ�W�;'��p����dW�/O�����}4��	\�`��O��c��t���ayo#���Pw|�D��0�?�u�_��12Uc#�a ��ݭ>����3�IyA��xf����������Z���n�@GPU n8	t��:��F��Pf�����@�N�;�'�=�,�p���>�5 "`��A��,������a�6��qj�GI�#Ӻ@��f*�5��3P4ဃ�8	t�:�����:��x	yo-ӴA��Α�$����*N�g�2�����u��>>KiRX�=�+���*�{(��W��L�J\�)<�{���ϓ���f��R����_�G!��r �0,F���A��F��g,��F�ڷsh�qq�6�����l5�ܴ�[�c��E�ms��׭�4Tf�5��-�����"�Z+��px1L�RY-G�}t8�F"��0zv̈ٟӡ�����#�C��[,��>��ϡl��[,��>��ϡl��[,��>��ϡl��[,��>��ϡl���vpm*7��xm�fB)*��t�e���g�Y�m�~e��="�Ǥ^�����0;���ϡl����޻d��l�|�(^=��nx�(Y���W{<4>��&�Tk�Q�?U��A�w�2�#�C���%]�f��'��d���C�B��d/C�@u97�+"��v:��O�p5��6���2<597�+g�Y��z���G�[���v�����_�dP�FO�d�FO�d�NY�吽NY�吽NY�����]�x����Y��<V�g�+a��x��(���+a��x���*���_������*���&�Ed�VE�d^���]�zk�/MvE�Ƚ5���"��d^���]�zk�/MvE�Ƚ5���"��d^�����zb�oLVM�ɽ1Y7�+&��dޘ����zb�oLVM�ɽ1Y7�+&��d߻}���g����j�KWd�Z�,���d����j�V��Ҷ�&��Y����h�����59TQ��j6pmG������2�D�4:�s��p<�nnnnnn�3���Ǘ�G�Dg�$��Y����`A0`�g<��(�2(��o�8&֔J�H�Iռ����N�X�C���z4b�;R^F����\�G�R_��}��ڒ�$��%f�r;/~s�g>�s�g>�s�g>�s�g>ԗ�$��+>IY�b�&)�J�BK���u��7��1�H��Vo\��k[��k�H��K�U�u#���Z��hY�g�+�H�BGwR;���������+�����w���n{Iz^�1��#���ƙ��/���͝\V���L��������/g��
nG��k<���}KaI�Հoq�v0U��&�ˇ�XWqtn|�6�m�{�ڀj_��������5��+>L�`�=�g8Y�����x:�����v]��>���>���>�P2ꁗT���<C��8�L��L�C��<Jd�c&�k/���d,�?t��:�������I��MɚU�v��)|7e�ᗵj�l�00>z��q�MI�VY	���%�7�_?N��WTo�cÅ9|9�ȣ>�9�^=f�p�e��|V�����(�d��c�^�����X�6���J��ov��t�ճ�KV�=��6Z��qT��O_ ܴ�~�8l�����9��M�����!��.�O�[z�K?Ն%����������c�s���0lan�De>��G��2�B��@ʃ�x	dӴ��	d�0�5n��f�O���v�N���"t��:���p�E���|F��f4��AӻN'I�$�&����I�MkNt��,r��Zv�^6��2�B��t/σ��:�J�Wg�W.�$�.��oǊA�+��H�� �e0q͎^�diC�pd�*�m"2_�d��K%JJ�@%	Oy����*f�A�W�K��Ggq}�J���E��T�tV�r����.����3D�Ǟ:5f�E��/�%�$��o�S�xm��RM��Rpm���t�Z�`��Ү��J����y�
��A�phx�e�B�gжY�-�}e�B�gжY�-�}:��C�t�r.�EӡȺt9N�"���^���X�����m��tg��"�Pd^���A�z�2oUM�ɽT7r�&��$P�Mܡɼ44A��t?΃'�Td�{?���e�.�H��k��:�r�'��2UM�Ȼ�<�O�S���8>�/A�B���NùA���6>����_���-���|���x5�g�Y��e���FM��z��)-�w({~��GZ��Kt��V�KKq����]����v�������^�_�k�z�|/o�{%�?�[��%�?��'�R��*T��!����H6���`�|lo��m�m����A��H6�I�� �}'��a���m�*�}s-��2�����̇'�d9=s!��O\�rܷ,��r�ܷ,��r�ܷ,��r�ܷ,��r�ݾO���~���}���a���~���}���a���~���}���a���~���|��� �|��ɿu�g�,��k�qZ��V�K[�y{}�/o����<����vM%��i-]�W1Y4S���Y4S�����2�B�C�9��?<���������������_�����>�bVI<E�A,�Vq3����&�&��
_2����T�('dJ!^�5ވ�"�jٝ���z1�9yyY�J�Kĳ��Ve�;/~)���j.������{��z�����$��%�I/�I�K�_��ԏ�~�%��Y�J��K�R?z�oT�덽{���f�v)�b�7g>6�u��\k^�kݭb�4�ٳ��ޤ~�\oR_[9/��1���{}/�j�����Ƕ�b��0��]��^����7�+���?�V���q�x����{߻�8�v݉�wquy%/�T����I�X��4Sgqo�Re�(,�:�ʱ}wv���d�%�욕��oʠ�������h�Ԏ�|���Q��K��ׁ���$lyǵ�e�v]��>���>���>�P2ꁗT���<Bbg��g13�u�P�4ɼ����ˣ��|��o���P�a~)��#�r��S�Q�ω����9z��Wh����~��n�n�,u�F����~iU���ҍ�&j8�8�uϱ��5c:ZdBZ�~x��O�V7���ۤ��U���a�R{)T��n��-��2ܫ�-���ۗ���Ӯ��T=�[O������~:30�T���gS��$�>�l�m������^c'��c%�0�x�>I�ئ�C��rT��G��o��qOV���GA�Y�t{X��Ƒ��+������t������Pc���|]g�Z�k�/%�^�g����5χ����i-��1셜t��_��9~8��IY1Y�C�K�{�/�Iߗ�$�mW�K{Jw����ጿ��ʀ��ޜ��H{Jv���\���F#�#���q����>��Y)�u��i$���^�)��e�5j藵	F����]���M|�u���^^�Z�J[��o�Y���͎]�+�q�8����ފiG!��H����`i&���J���{J�g�h9:z�"�Td�
��C�t�r.�EӡȺt9N�"���^��A�xh2oM�ɼ47��&��d�:�������_:���S��PdRZ�����9gr�'�T��ʜ��S��*r~�NOܨ���5�*��a��|�v�V�����[�NE�n�5>�1n����=�<^+c������쟡o��m�o}vM�ȫ��������}'��I����1�Z�c%�v�}��C��d9</Aϕ���)+�Tl/o��Hq0��Y��p=P����)�5�*7�-�tt�����[���q����!��d:OL�I��=2'�[��Kv>�U���a۬`�u���iQ�̇\�k�o�s-��d8��[�\�q5̇\�q5̇\�q�̇���r�lo��m����c+iV2��a+iV2��a+iV2��a+iV2Z�_%�;	-J������W�i�KR�䴇a%�:I-!�Ii�KHt�ZC���$���$��I\�v5̷c\�v5̷c\�v5̷c\�v5̷c���~���|��o����+��s]��b������q�����t��I��t���_���k��s]����-o���3�d��������'4'7ޯ�_z��Q�(��"O��, �ȕ|JY��W�NO|�&�<�dMd��
_2��$�@�H:�WkQM�WM���z1�}��s�%�LWz�w��p	����~s���+=�s���^��jG�R?z��ԏޤ~�#���H��٫�j�֫�kٱ]�ٿ[6�f���͛��H��G��ż�_��Q�67s���]���R��6��ֳ�C�$��������ke�������������S�Z��(��Ww�K����/\l���cj�����6�ݻ{"��099B�yY�ke*��_��M����y�v]j;Hd����Ya�u��<F������Ѭ��59�;?���}�Y���oU/W��Z��L9��GK#D���Y���x����x��,ˡf]2�Y�t��K�x���bg13�rw�9;�M���&�+/'Y���n�����X��ۈ1�g+�q��?U�w��i|ɮ՗ã�]�ty���[�tME�b�Ye�đ��:wO��!�fͣ4j��U�K���^��Jݱ�$��@�Wk�U��&�Ҭ��ܛ�-���ܟ�-������vM��{+��ȭ��]���z���rr�=�.��V�+��yѕ�����OzG�{�����CO�)��NqZ�$��M%�/Q��,��e(���@��\��[܃zr[���h1��x�м��B����W��x�_����_��<	Y��������TO�r�w��;���[�z?|���G;�����p`?|���T/-x{����g;��x���$�K\H���7��js�������?+� �t�T����{�WX��W���Y#�\e��l������o���A�yM��,���F�o�z�O��9�a<��Ah�JA��z�k��6���Y�X�qߎ�٪��I[S�p`�we���`Db�(�:�Q�J�IW�=��g��y�Q�t*2~�FO�� :���� :���� :���� :���S���rUNO���U9?��'�T�������~�P^������d����V�<���'r�a܊��"�=ȭ�r+c܊��"�0�N7�S���c=�X�dV2�����>*�L���x2O���k���
�[�~�:O܇	ܨ�{%�(^C��R�{��OM*�V�v�a��v�[����l���tq[+a-��_%��Ύ;c�5|T�[J��d8�6�湧��2ݏ�!�t���L{����$��2KR��
��+I��AziP^�tO���D�m�>�tO���Fx�Q�+to�;��zc��m>6���IiKK䴷�KK䴇	%���ZC���$������Z�%�8I-J��d8��C��d8Ύ;��bz8�oG��㱽v'����q؞^�I�ۣ9{u'/n���Ԝ��3��Rr���[J���d���%l�+d8�[!�J�2V�q�Z[����l���d��%���--��in6KKq�̇\�q��*6V�q��C����L���el����}��_x�Wގ��Ңyy3���yy3���9y3���9y3�g\ι�:<�nnn�М�z��}ꂁF@�|���>���($�	_9<��+�o��}|�<M�x��Q��F_�HׂP$I+m��n�z�qM�8?v�׺�=	/�g>Ԭ�1]�K���r_g|�����{��cb���s����?+�?z��ԏޤ~�#���H��G�X�͊�߭kݭW�q�W7�f�l[͋��H���_e|1��类s�ݮ68d�����%�w�5�`��5-�>��ס#�Ow�t���~�S[�)��S��[�T�N�kc	!��r�a��;ͥ�ƶuƶ{]�y�C�U��V�d>�r��,��f��q�Rb)�HS�_�@ǳ�!)[/�޳��A�%~Z������7����s��p����]2'ݓ��mv)��VwUQj{n3��<W[��)<z�Y���˼}C��<}Beг.��t,˺]C�� �&pc81���������d��rs���Yx�Y���n�����F���,��P�[�B��.:�q��`���H,��d�������8q��/�]��������#��M+J�X�2F��_���v��ڪ���!k�8M�e~Kr�V��8|^��Ƚ�7�C���r���E�ɽ����"��d�N��S���z^���߹���qZ)L����En�9�V^��j����*<�g�s�п[��P�5�Z@~�R��ۼ���4^oq��̣%�x��FF������o����@t.NI���qҷ����,㤴���|��`Ď�|	���V�%o��}9[��<~V�8�K��p?+zp
TMs+}_�-�n_����g�q��1������8�R�A��0})n��l�7����#��S�ke9����jV�?	iFn��}�n�����ȏo���"S�j$��˿��� ��e ��bjѸ��v�����h���I�����lW+�ҫ�q�����׍W�}Ƅ��z'2�$J�B�ܡC�84<]E(ǰ}q��NO�J�q쏜{#�C��Pd_:����uUF��S���rUNO���U9?��'�T��8��+_�����8��+_�����8�}sZ���2��V��]����9zg_d���{뱞��g����{뱞��g�+��x���(�����-�x��H6�	\��:Z�?dRϹ Үb�i-!�tt���wD/S����iP���
���ktg�n��iT�=*�Hv0bC��$:���'���n:�"��81�B�"����õ�u�d-����}k���x���p��Hގ;+i_��ι��Ikw��w��;��������|�㰟��'���AziP^�T��c�Plv
KGa+�̭����̭����̭����̭�����2���Vҿ��W�-!�IiKHp�Z���~��߼|w����~��߼|w���۠�;tGn����]���Atv�.���Ңyy��D��/J���8.^���pR�C����L���%l�+d8�[-���2V�q���+m�R��+m�z:Wގ������?<}��n��Ҽ����}+�GJ���Q=*'��D�t��>��۠��@����	�	�	p���q�gI��O��X�N�rxE�##�"&��ڶq�d�j�y��z�?��7ȣR�D���bۯJ\OE�O�a��sE5�~5��{Y�N���֫��덥�e/\l��[9��o���ٿ[7�f�l߭���~�o���ٿ[7�f�l��͜�خ��֩z�1��1��G�n����vU�e����;eG8���l���S�wmJ̈́'��v�iy�Ywy�os[2�^��� �5i8���W'Il�W�$<�n�7i����$U�E��!"�����q\��%"���Σ�є�K�1b���/]�d�����q����V%�X���oϣ;a����E���DB����c�z:ǳ��q||�H���G�a�[Z��&���wX�vx���c����K�a�=dv^�.���.���.���.���Y�t���M�|�_5�y�̺��h�����e�����9;�y_�$a��7��G�$$�%��/�Ԩ��O��`e�˯�F�>�����'�ß=4*
�����'�ٹ��t��e;}^�FM��@�U�^�:�:.��=�wd�z�D,��lz%���;I�������G�A��Wpt�>�vσ҈�3�t<��Ϸ��ɥ֦�ȥ���o5eZ�d�F\~��)O��t��Gy���56M�V-�ee~6vS�r{Z̅UΎ�!�0�����~��O�-G8=��?9O��z�yk�܎@p������T�$w��<=��+:9#�	����V�o�Ee��4�?������������帬���)+`�@���[�+d���R�x���-�:��5Og[�g4���[-R���^��bm�H����7��l6p�TSi@���X���/a+��'Բy|��&�7p�1�K�As����X�}Ǧ���>W�R�xiy�^��)Y[.�LMMmԫ��L���?��f�r٫(�3�t<���l�����z��C�x�2oeY����:OU3�A��Ec}��O}v��]���񰽾6������^���a{|l/o���񰽾6���������}�Kq��n�J���|�����T'�;��y���R�'����-�x��OL������>�U�J��m�?�UĖ����?��R������	�����wZ敎���Ii���s�k]yzgXYY�#�}k�O_�^Ge"|	n�G��qY"O+n}��+W����;ae>��C���V><�ֹ���2�����d?<�v�P{*�*�kV0b����-t��u;������Z�q%��Z�q%��Z�q%��Z��KV��j�Y-Z�%�]d�k���y���x��81O�)���?���pb��S���ێ>;q��n8������|v㏧����b��S���X1O�)�`�?����c�>v����1�;��`|����c�>v����c�>w����c���n����x�t'n��ۡ8�w�>�	�ۡ9x�'/��㰜���/n��Ҡx�T!�x6����n���`|W��	�Ҿ�����P+P5�P+P0<�n�М�nnz��Q�g�t�������$�a''�k�a썗Ȃ�"���폛��n��]���ԛ�	�H�`�F�/|�e��;v��s�����}�y�~���u�޿Z��g?�ҏ�i/��K��s�l߭���~�o���ٿ[7�f�l߭���~�o���٫��9ٱ]���T�����������{v�����u��:�9Ʒ7���C��ke��޼mo=�έKe}K[������A[9Ui{Fq�Ǽ���HM�=G�3���jsH�F�]��v��h�'(a���YUGc/!��8�������f�e��z,��i"��ҵ�5��n�E��B�,���;,��c=�X,L�a����IY�=���FT���m��d��[��,0�L�a;g�R�6���6uv�P}��^���Q�6�r���w��x�w��x�w��x�t,˺]D�&����j/�����f]%�ٹz}�)�YA�L�����/+i���%�/��[�Ii��h�rxb�lДWf�_�i�fjƲ��m�i1�����mv��]�ХQ��43Qph1?+o���Q���;�g<y��k����ee*P���l��t�|{o�A݀�΅��S��Ws�z������ɺu���r�[+�N��H��
W��iD���	4jⵝ��dvZ��"4�Lsk��A�P�J��x�&s��V��Lo���l��ܮ#
&�Q�x<G:_g��B��b>�6Z���߹[���=��9�x>w��Cǁ��>�W��+�|o\+�+����~pc��B���H�^GI��%n)���Ĭ����ޟ��B��"�O��t*�����no��m�D�*����[��=r^���l�0|G���؛~�/�
��4��=����B��˿!��b��d���xT�e ��`���F��;���㸄�//���þQͯ*S�b�5*߮�!{�2�|SS�\�]�Y]�1(�z���Ty%��A��Pe]
����*8���S�zj2M��A��Pc}��^���Q����0��&������d���RO�C���=���[��Kp^�n3�-�{%��d���9�1ްm��J�\�z���9-O��m��mk����m��t���*��!�m��V�敆��a�c�����;�K[�r��\�*�����1Z�$�|}kGO���j���<}*׃�+k\��g_F�++08�N����e��q#�R,�����gގM�r�*���2<����G>���ǒ0��9/����RH���`�S7�L���(�4�>kGZ��ְ�u�=�k��a��]�k��-trE������f�険:fn�����3x�^k�Z��V���^jׁZ��V�x4�~?��O�����4�~?��O������~w7�O��Gsx�~w7�O��Gsx�~w7�O��Gsx�~w7�O��S���~?��Z��)��
�ǁO��V�<
81O�#�b��Gn �?���A�X1O��������}?����}�D�h��w7���S����ǁ�-�0b;�G��G^�H���zY#�ޯ�_z��Q�(�3��8�3�������������|�o��g挲���d�j� ���(��2#W+D�굴?%/l�h�l������nn7�cƱK�8��Z�k^�kݭq��6��ָ�׻Z�l߭���~�o���ٿ[7�f�l߭���~�o���٫��9ر]���|o[]��]����^6����j�o2��͕��SW�e/J�h��tH�t���a�����,��yd;g	����=�?g/Q���jz�;����~��"�I���mo}�������v�G�#�����]�����*{;T=f>6����I�9�*�O#b3Yk	K/٩��҆�;��ku���wc�Y���ޏ�Z�%K�+��N�gd�콜S��߭�]�K�7�w����N类��K��=8E_�?a�p9w�x�w��x�w��x�w��t���M�K��,ˡf]�ֱ��D��������M����dj���/��^�d��ĭĿyG��W���õ�p`Q8V9�*F[�^�����=x^���z��0��/۞�m멥����om�=j�z���5h�(���wVU۟�J^�R��8��r��9<U/FYӠɡx������}U�>�FEШ�x�=�^��S�9�`8��܋��Q�pf/�k�fVS��N�?--T���J��%	N������W/%張�6j.���M}�m�v�>�q�[��{�Ϝ3���^�E��P��-����r��,J�-(�j�9��Ř�{�-�pb���W<�NV��G>x����m����1+3����`�1>u̖�~�|[�����C��z�M�H5�6�R�F��@5^�+��mv��K+��`?v&C�[zˮݻ�E�tvq}zԥ�A��;���)�9Gݔ��=�%�6�A���j_�ڰ)|�����9{\��yx���s�G!ո�:-C᰼z/��/�RP��2�o�q�G@��t���������x��S��T�Ȭ��S��jv0mN7�S����`ڜ'����S����Kp�)n�!����4�H6����i^q�?�t�;��n���|���?��ݺ��Z�d�]?�GO�����3�a�����3�%��>�k����i�|�>H�����j}�^�W��0�rE��������i�j2p��}@�Q�5Z�#U�K�Đ�C��]�i�|"��f��k�#y����>���vu��肮+Y��6K����-o�BA�d��dx��Y���Vsx�F9��#�p�F��^����n�~S�L��S'#��)>�)>�)>�)>�F���'���zY�K#]�dk�-f�KY���h���=-f�KY���*��ʽ-2�KL���*��ʽ-2_��K��^jׁZ��V�xFoH��I�	#4,�0��Լ,�0��Լ,�0��Լ,�0��ԿKZ�������]-?KZ�������]-j�KZ��֭t�Fn��k��3t��],����Z�d��-j�K$f�kV�Y#7KZ����Y#7�L��S4x�����3x�]-j�KO�+R�/+V�ej�KO����t��}-k�,�\B�e�,�\B�e�
'��|�'��?�I��O���]�����������|��,�}%�O��7��j�AQ����J���Q�SM��V/�Jj9�0��X>��Kb��g�����Η���c�[W�Z�ln�s�k\mꗽR��_u�����f�l߭���~�o���ٿ[7�f�l߭���~�o��\l���\lԽk�z��o��o�oj�wjò����/i�K�tmrJ����镟��n?��E2�q!֠�5�ek^+�Ϡ�����t�3�c���;v^�J�����,�<��&J��7�<�v����AGv-�w6'cq$wtH~�u?E���^粣��U���)���~�2?@S�9Æ���l���씳ۨ�{d�n.���n�f��7�kko۩����v����n���6�~­�/F)�;g|?g/���|�p?)xY�q����p�q��q��x�wK��@��P17����̻��<����������k/��dj<�R�/Y�$_����Lx���yI��4�4'v����-�y�z͇�g��|Rh�k�-�zS�!�5�m�{��=?���֩9��o�Ы�_G:�O�Z�u+M�Pl���)��?���^��S��d9!�B��UO#�A���;q\N�+����t4�G狆�D��	HK�����$ⵞ�?�����Wz�(G.r��R��2?a#���Ll�R(�<��1����]���U��Ky=��s��������C�◜T��,R���u�b�-�"�:�o�[��:��J��5{~��n��+�5f���Wm��u���E$�/8��8�^ql�H�}yA���>Vbk4=N[Q)V�|���v�d�t�O��R�|b<>턇����]�v6�r���`{a���KnG�|�?���d�� 8���J��"�09����i��̾r�-��I^�d~Z�o�c�/{������T:/��=T=��z���z��ov��o���l=���7�-�zm�U;����m�v���_ݿ�s-�W2���q��\W1޵ͻ�s�%��$�>�KGtJ��9[O�+k\�m?4��s���Ҷ��V��t��>R_��c�d�Pb���H�|���%�R��L��S*��"^V��EځL���<c��<��bF�$j�F�P)��
d�d���2Vo����f��YT���8	!�S)G��Z��k��F�+$h,�F��q11M4�R��i��$m/��%.�
�m���)��[��_/2?��d�⺉z�)�9���;�>&9���k<�nSG$Q��R��W���z�Ǭ�z�Ǭ�z�Ǭ�z������������������o��7����y�#]��k�<�wǑ���5�F����zZd�KL��i��-2_��Z�r��\����/�e*���<u2�L��S(���<u2�L��S(���<u2�L��S(���<u2�L��e*��J�vR����e*��J�vR����e*��J�vR����e*��J�vR���$l0��jH�ad��e*��J�u2�L���.�9K�R����S-q��\vS����9��N~>S�����q�gI��O���N�v�������$�>�>��g,�9g�ɠ��������<$�%��oش�o�}-�R�펎7w7{Wy�q�-�ɼ�6�&�d��ͥ�������l��s�k\m��q��7���[��Z�k_�k��~��ֵ�ֿZ��Z�k_�k��~��ֵ\kX��\kT�j��C�����{ڱOEX�w��j����m0�t�~55k�ی�˟wa�c�����Kv4�V�O��H�T��|{[�=�W���{s�5���BA���u��eR��'��1ie6��S���l���Z5�V���OcF����݆5�������T�W��[e�n}b/���ՠr�-�\�N����ˁ�笏��������F�J�N�I�
��[�ծ�R��r�K�ܾ8~��/�}K�:����ч��Ê|���'�������������ퟏ������r�z\�ޗ/vl/㽳�2r�W�����]e��Ӄ���FV�t��*��Z{)�^;:�KY��՟�ujO��dޚ�����n��=V����[��{�S��Q���ᕵ�yźÕ��D�i|iѿe[R�9��#d�_�+es�o�z��~w)t
�߃�ʻ�݄���>G���%�ھ=��K�y^����X�c���|l��_F��Q:+�fVI�k=~#��%t*RWB璖�ظ�-��|�t��������II�_n�ҳ���ǁ���$���*C����)\��:��;��s�Mq�zj\n>K�`������������R�7�XY%�/�p���b��G#��6T����|���BA�8��S����BK�lV+���$o��|�F/���@w<Gze�C�/W�-졽e�nݰ���L��X<��_���oСe�ɊT�2����9C��3��F�r���yK�aǛ�E����+����:�K� ׅ�y:�/o�Il�O���q���r[��K}�����!��i^t��܇��s�ұ��X�t�uͺԖ�f���Ҷ;�V��r��\�k/O����:��H��ְ�9I�W��K�4ʾR_��U�r��R^d��	�$f�d��R�KY�P$j�R^�H�|���L�$��V�e(����.M�H���2w�MXY���d��՛�����Fx�9��9��9����YgFs#1I�����e�잎'#�?�vN���#�R59�����e��"���?x����qm}`�0��Vb~�>V����qC��d���S�)���r�|C����\ⵇ8�ρ��ˁ����������������N�'���������rs�rs�rs�rs�rs�rs�rw�9;����:�w����ux�^;'W����7s����fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�fy�f|�#_�H��5��#_�H����N����d��:�f�Y��H��5��fx�fx�N��vGVj���\RF��+8s��lⳛ8���+9�|Γ�����}�$�a'a	;I�BN�vU�S�}�����Wɢg�<�J%�'H:�B�M6�wj��K���we�[۰���j�ޤ~�u����y�mvJ^�K�6�/[:^��޸�׻z�w_����~��ֵ�ֿZ��Z�k_�k��~��ֵ�ֿZ��Z�k_�k��W��Z�k\mjG��5����j*��e��[�����zf+����H���L�bb~X��	#�&[��ۻ6G'��
�������^��n��Sa�r��Kt��Y���u��P�`�Q��H2�nJJ������m��ųi����ݿ9���}�q_E�]�[g+������7o�:WKs��N���{<����p;0p�i��=Dg[:W�'坄�ӥ�FE��I�\G�<������8v���//��(⺉~7��;{F����3�k8���k8���k8���k��8���ώ��l/�r�z\��Y��������l(���0c?���.>FA�pbF���Q�kW��Oe=짼U�sZ���U�+4`čW��U��e��_v�z�w�A��t�3��h��[�l���S�k���E���u�_4�4�߆�^_����4Ck��[�+>6SW��v���~�_�!�<V��Y�g��2�-�x�G���.���������iK,"������d���V��e�q��Dk�L ��p�K������.Z��xi{I!�*���x2hoe�a��è~�w�Z����sn�J��8�����^qC��0�_�s�xwA�p�)��܇���������LW��\�V��Pb�ƅ�*_��<	+$���}2_���~�%�L��_��\b�o�G�t:q�C�un^Iim�T��8��Ӷ[zK/����k"To����)u�,CSr�|�.L�*M ���d�+��Vv�ۉ}su�	k�h*���Z���T�]����=U^�VEܩ�=�:��gжY��2�M$ë�ް�+��C���h�ұ�kvi-�+c�k�}X6;F�уc�u�2Z�W��K�t�<}3$K�4ʾ2��L�2�`�R��Q�$k��w����5�F��H�|	�#]�$k�v��,���2������/��h�̝^��F�H�|������)�j�VVo��s�.�&�q(Y�����e��z8�&x�M�d�M�b\%�b\%�VX���riY�p:������g��;/q+2�s�G^F��l��)ͥ6z��MO)�#�1�ݑ�f��Xj[O���'�	%�T��NY�D��v���x�K�J�BK�����5�Yp99�99�99�99�99�99�9;���N�'���������5�P�5�P�5�P�5�P�13�13�5xE�Qw��]�5xE�S<S&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�2lS&�5qME�SQw�]�13�13��4�ɥf%+1)�����9�ݕ�:2�'FVbj�<x�O)�Ǌd���F�F�RX�XBN�v������}����g&��M;8�cV�À��4�D��)���{|����_�ݿ��{��6�og#�d��_�ծ63�l��kk�A�k��K�~���o_�k��W5q�~��v��ֽ�׻Z�k^�kݭ{��v��ֽ�׻Z�k^�k��W��Z�k_��Vl��;�;�d?m[tV���WmѴ�����+=��)L�-�x�W��Sq#V�14�~�k�i��>%-���Oc�[���eP�v=����l��u�M�c�r���廻��V&P�)[��D����6s㷩�b����+���yo-�Yݒ�;�(�l�'r>���x:�l���٫#r�QY�Ô�d��>U�/M�'�����a���/[	A�Q��a1\O��/2v�S6+�����ݢ�b������k8���k8���k��8���8�l�}��/w��݅��l��_��n��L�<����|��+*�Yq�E�~Q\�Mi�̌�i�6;F��A�������6�����2��/���[�����:���U�+d8��^��9��}\6�V^�F���셯�Q�����-�J�����\��Z�_�W��2/]��Z���/S�}�ft��UحUg�gM����jβR�Q���������j;�̗�)(|��T�w��>R��^C�ʮ�IJEX�m�<iY��J>�����J�+h^<���}Qo�q��{���=��R�,�������x�<�����+#�~������OG��`ǃЕ�lGy\q�Ď���ߜTV)���t,�b�/��,��;�_�`�~���3�Y+�ՙ+��{�t��ЏV�U-�+Sۢ����Z�����FǶU��ie{e������z�ׁ��n%�%�y���l8�с�W�?�)Q�A�n���*8>�}����l}��d/-�z��>�W_L�W�O��U�Ү���[n�������[OIj��Zzd��Hzi��dk�l�G���9F��H��$i�
ʠVU��rn�&�rn�&�rn�&�rn�&�rn�'<S��6xE^QW8�]�=�����=f_Ǭ����F��d����vq�x����p9{�mYY헕�
��Q|��3�BVj�P��v)�J�BVj�%#�)/�p��Q��,2�њK�9�}n�SQ����|�B~ݗ�v&�+��|{c*Z�Hv�����f���=����55-�Ĭ�K��׃�x�s�~�����Ĥv%#�	�H�BGj;P�ڄ���#�����;/|���#������]�eئ]�eئ]�eئ]�eئ]�eئ�x��x��x��x��x��x�&x�&x�&x�&x�&x�&x�&x�&r;P�ڄ��$v�#�	�H�BGj;�ؔ�Ĥv%#�)�H�JGbR;�ؔ�Ĥv%#�)�H�JGbR;/|���#�����P����ĥf%�������ĳ�M��w9���ud�'��Z���R_Qj7�7�7�7������v?VR�%��F3�]��VB�l��esP��0�no���d�l���#���z�6m���ֿ[۲?gF��ݮ63�������a=������w^����W5q��q���f�k^�kݭ{��v��ֽ�׻Z�k^�kݭ{��v��ֽ���Z�k^�k��I}��?gFݫ�U��٥e@�Է��ݍ��ǭ�;/O��{;P|�ڞ���ю[��HyL��?�/���?���igy\��y|��\��P�W�{�z��!���g#H5,V�$[�,F�7S�͔�a�op�;��+6-���#�J5=��"P���4�*ŏ*�K�OFĤ+ݙyJ��ő����߷�$ލ��C��5�H�F�E�I�}?>ݍ���&6Gd೏��#\t�Dq����g$k=k��H�k��O��O��O8�NG|��z.������������5.���}������5�#O����VU��+/&��)-LW23�ĥme��ݨtn�����S��]��j�H�ܷ��D�c�Lx���ꮺۣ�\l!�?�Ns��陼�ڲ��ܰs��~�a��6�Η��ǿ$��������^���u�՞)���$n.�����gN��ԏ���V??8l�}���_����~s]��!4A��O���Tq~���J8��Z�b�I
���Yć)k�2���VD��KJ�!Ǹ����9>pĎ�q����zx�K�%gG��`�q�W>��KE �=�E!��%�D?a����HV�#�9o���Ti�/�%�mvيǾ8
�1)u�R� �?�����,;�P$w���H�܏�p�����2V/���]�Ȧw�Q�@u>�U�?�l��nר�hNr>�$t�~�?�(nX�h-��L���Hв)��V�<滆�z�f����|�K�5��9+�����z^ʍ����a>u�Z��KS-B��H�+rn�N�������u+i�>���N�HJ�!�m1�ZFIj���������P+7����K��K��,ġf%1.�'>�&�rs�rs�rs��s��7�����+=S�~)�Vwo�{��wo�=ef�Ԭ�a�5s�E\�aw�NK���ɜbYơ+2�d~�_ݰ���a��
�_/v���j��1_j��1_jK������?Z�s�g)��E/���u��]�m榌�����yԱ0��e�Siq��c�bk��r_QIK��H��jA��������wi/ �c�{e�^���������a9/�g;s�g>�s�g>�s�g>�s�s�s�s�s�s�s�s�s�g;s�g;s�g>�s�g>�s�g>�s�g>�s�s�g?)�>�)��#�7qME����j.��M�SQvGbn���Q|���+5���Q|���+5��BVj;P�����%f�#�	Y�H�BVj;P�����%f�#�	Y�J�E�Q|��ݕ���f��/��Vj_�r�WP���侢�/��9���us�E/��%����ԗ�Z��FA# �_Q0H�$o�$�ԓ��dX�,2d~T���ے����Q�lj�l����v��������1�C�q�C�1�C�1�C������l������޷���f�l�͛y�o6hcb�6(cb�7��7��7��7��7��7��7��7��k^�kݭ{��v��ֽ�׻Z�k_�k��q�s�ln��4x�;����5F�a��1u�K+��$l�a��]���j�ʝOcF�l��}�ܦFW)�(V���o5���ߴ���P�b_V�ܐ�͔v�ۉ�S`���-����䭗<�U��a��)y/�� �#���\���̇����i2x��,62
5��Sv��{}~�Y���&�����lw��kt�r��p)R6��i���Vv���}�&�e���Z����@�62�=f�=fYS�BR�����f�\m�O>_Q����Vwo�r�mc����q0=.�ԗ�=ކ���j�P�2�a>/��x��K�t��K�t����2�?(��-#$����?(���x�Bb^*}^�?����L�%�w`�"�HA�C�JJ��GP���d�ϕO̫j]v��y�.ڵ��E*�ѕ����r�<�r�2�,V�
�jd��FR��lx�����%eCzsz\�K�����k�eU�^�e�/���U%�ѱ��C�Ӿu/Gr�)xj5�Uv/��}U�o�� Ś�J��dv�%c�V!rҔ�,>\T�г�=8�,�{���缨Ď��5̣%�N)�����/���/w����}G�e��V�#府1n�����@5����-�vYn�\I.+��>7K���<1*^�C��8?���ZK��U�[����+��}���e^�W�$m�����o����=gn9�]d}��e�P�.F���^��7�,�i��O�4�kx��_+�����|ӫ.�̗�7�O�����ǧ��1߲�;����[����]��k�d���G�$_�m1\��Q��}1�����d���:�����M���1.;Q<S.�2�Sa>a>a>a>;`���v`�6/~q���l%�L���f�5x�Y�g>�;]�)�����)/Z��z0����?+�����]�r�=���|e������SQq#��jy�/�ݗA���]��$���;a���R���\|�Ϣԗ���>�;�l�C,~흮7��ϻ����L�Q�J�����G�C�y��I��>�߈��wg#��B�b����m�?��|�?Б������vr?�9ݜ���G�g#���������vr?�9ݜ���G�g#�	�b�&+�Il俶r_�9/�+�b�&+�b�&+��1_E��Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ���Ɋ����%������l��r_�9휗��G�g#���������휏�����������q�C�1�C�1�C�1��_\{j�ڵǶ�q��I��XF,bT�KE��}�nL��[m�^��/w;����q�/v�o_���]���1�C�1�C�1�C�1�C�1�C������������������v��ֽ�׻Z�k^�kݭC������������������v��ֽ�׻Z�k^�kݭ{��v��ָ�9��4[J5���g8wv����V)�o�����-��6Cη��5<����C���põ8j[�#'&��<�vDn�����孰27��[c �,rx�J~&ϕ�ݭHx�*�&��l����e�VC���t[���Y+[L�gI��D�m��{-Mn3__5�l�X)-���W�d���?#V%g'+S�N�X���P랛i��H��϶U���gr�^��NO%�+��������J�Kyz�n�g!��$=D+�#]�l�wv�s�H����oKO������u�}�^�������e����{\�|�|�|����>]��'��N���k/���.����/���|"�>H��L��P�jN�'��x��{�����[s��Ϲ�5[�R�3^��AGFo���-]�ܾ�2�/���q��.'Y"�X���x�~YWy����� ~�e�W�������wc�������v�Uso�k!��f�4��8�����0�v?�� 8�C�C�ž�F)����9/�kqy���K�=�yY�J�����}��|o*?k(0��Ix<13��#�~s��?R����%g��l��k�D�K�R��4w�'Z���ME2O��0	Y!�P?�B��);�?C���/+eg��K�8�:�KqYA���/v+��Y��@t*�m���}k����v��;�(D?�X�Խ[��4쌗e'v�r���x��C�-�$(VG�<�%W��;��m-@�я���j.X�39������+�:�[����%l�FV�t��4����Q%�g/�x23���e2o��4�Πbg1.;�1,�P��t��O�ߊ{o�=������w�|ɜ{Yǵ#��軜�(��D�s���ɜ�R?f���0���/��ɱYk��R���l��n����������\|�����n HI��\|�ý��G�-q�k��m�����W?j��mw��ke��<{͏\W{	ln!���ci|1�mu�nzڴ=n8�Fq�������ʍ>2K�|P�슃��G�0���#��v%ˡ�m�?cV�ޡ��G�g#������?{|���#������?{}q��q��q��q��q��q��q��1���Z�k^�jޡ���ݟ�?�v���]�����wg����ݟ�?�v���]�����wg����ݟ�?�v���]�����wg����ݟ�?�v���]�����wg����ݟ�?�vuǢ���}q辸�_\z/�=���E��m�׶���w������{n���^۰���c�|1��_|��>W�+Ꮥ����ʏ��G��I;�
O��ݯv١�LB�v�<��:V���ҏ�v�aV�K�u�v�o_���]�����wgoP��oP��oP��oP��oP��p��p��p��p��p��p��p��~�kݭ{��v��ֽ�׻Z�k^�kݭ{��v��ֽ�׻Z�k[͛y�o6m�ͼٷ�6�f�l�͛y�C�h��+��e|��$��\|��l�a򍑤>Om3o{译�6�.�/D��g�Ȳ{y9*���)����nTl����p搩���-'�2P��er��-�]L�wM���A�ݕP��v1\��{ip�+����t�
��e����K/�צR��*�o�\��0%^d
�'��׳+V'�^�m�����6�&��S�rhn�g�vF��H�+�������6��-��K�z3C�T�?D+�	���e;�!�*0��ݟ�b�������pG�F��>]dv��+���f�kR?�<S{w8���%g��|��{Yǵ�l'�{g�l.�}.���.%�b^%�b^%��%��c.���[YA�u_ߚ�S'�֯�V�Z���G�$_�%��d��TZ��QK��z��q14�usZ��\5��m��A�ܡZ��ZX�\�����/䏡�}�d����-[���,1}�(VS���V?Ӡ�z8샴�`u�	*��s�D ڍ7�n���v����r+�����%�c�D=���&&E�V�]�x��s��?R���$w�G�o�VW2?�eg�G\H���VW;�W��R�y;����4��z�[!�:�Q�Vd�v��]�e�u�T������̖�z_����W��1^_����z�g���x
�GI�y��늁��b���+M����u�/U����dt�Gm�M�u�l�+�v�e�4<�/{�qF�%�:�&Rۭr���g^z'�	�
�;�yy{�y�՝7�&�ߑլ��))�w������OIi!��/�r��ܤ뜣�����k*�YT
�d�.%��].���.�~>]�����eئ�yϵ��Y��y����]��)�)��q�H�jV|����w��w��ڵ�΍/d�}�7�d��ۿ�n8c'�GWp)u�(ww4?e=��#����m��l\w��oX��:2ߢ����s���� �:�(���)��#��`��/{V�Aq���%Kb��T��۞ʍ�i/������0��4[�b�6*^ƌcj������6Wԫ�,V��S�Xֶ��~��[w��C���B��Q�vR����׻Z�l����ݳ��g?v�~���9���m�ƶ�c[|1����ko�7��lT����mvm�͵ٸ��Z�og���y���{=��{������7��og���y���{=��{������7��og���y���{=��{������7��w[��y�o;��u����z'��O�蟻�?w�~�D�މ���z'��O�蟻�?w�~�D�މ���z'��O�蟻�?w�~�D�މ���=a�E�c�v�]�@��Rn����bJ�O/[����4@66��ڻ_��7���)}�/f�oP����θ�_\z/�=����7�v��ֽ�׻Z�k^�kݭ{��v��ֽ�׻Z�k^�kݭ{��c{8c{8c{8c{8c{8c{8c{8c{=�ͼٷ�6�f�l�͛y�o6m�ͼٷ�6�f�l�͛y�o6-�ż�_��$���Yʻ#�W�$��+�m�]e�<�8m��$B_M���z)#�+�v���Zչ�7�ԩU?Qo��e9_�&��B�y��G��lC+� �+tݎ�')�e���;=Z����B��������b�\0���d�ŋ��vt�.�Q�M�H�3����X�l�E@�߅`Ye�G�</
��Y�b�i*��B�m�*�l�{�����j!Yk}o+Z�����?m�+�����)����y�c�y)�J��\�T[J4Rݗ�2��f��s����ݩm'K�_%���~�qʜ1�~�s�5��͍��%�����s����wu�z���zw�~>���>���.���>���>]���u���̑w����iZ+��ޗG���H���9��s����{"��\]����uGZ��tD��{;(�����Z��+o�U�V�Y&�}VR�i�)KW>/
���j�k�l7"�G���;}�>�Z�lb�I���6���-J����8��/$J�\����J�Y#�Պ~�WY�դ�ϱ��C��n7Ƒ�q#��Y\��^�Ď���8��);�Ď��Ǧ��߸��C��?�k�����8��[��5j!�}Կw��B���}��s%��W��Iy[\g2[9�=2;��g9�K��/�P!z���2;�-�`�:d��*��gb-2B�u�Plw���g�	#�+���U��G5K����o��!A�t�#V%X�[7�#�;m�ݳ��F]>i8e�a�V��y��S���wGA��c�~��	��e�c��}12��)8Y#<	��Η&�q(Y�x���pw�p�����8�O8�O8�NVz���{�W��{��{��w��w��w��{�Y�g=�s�H��ٿ[9�+�ͥݮ���ak9�Q�������ݹ�p�q?a���U~�lX����g:^�|m��ъlR;��F���ݳ�S�����;����^6�̬��k��:��6ٲ���K�yS�lhԶ2��M��UXv�������W�+�CEK��e��t�v������������V�6H�vl�5=�[��sީ{6+����j�����[]�y�o6-�żط��b�l[͋y�o6-�żط��b��P}��R�*^ŵٶ�6�f���mk��q��6��ָ��Z�k\mk��q��6��ָ��Z�k\mk��q��6��ָ��Z�k\mk��q��6��ָ��Z�o\mk��q��6��ָ��Z�o[������{=�u���y�o7��w[������{=�u���y�o7��og���y���{=��|Q�K_)v;���J�?cq\e�`�$1�H��K�X��\|����֡���ݾ��]�=k�E��v�c{?v��ֽ�׻Z�k^�kݭ{��v��ֽ�׻Z�k^�kݭ{��v��ֽ�׻Z�k^�kݭ{��v���8�Gh�mm���q��6���8�Gh�mm���q��6�K�_��_\r����/�yS�vHch�i�M�?�#6��M"[i�{�Ken��7?-��-�G���������64���O+,�{y�W�5���oSg��v��g?k���"����NA�u�1�^vF��~\91����[��%RWl7/ ֤~S{A��B�]��V���$F#����eנly#��V��JB��zl�w�����+��[�I[�}��.��ݕIZo���g�Y�b�[�Z�ʻ[�6���)������Ӝ[�)���y�팽q�o16���U�l���Tw�����o�l��*��*����ث��ٱ]�K�R_Z���)�p��p��p?'�p�s����c�r����h���|W���W��D�=�|���+)ZPzV��������3���z�uF��]���&f�f�v�۩�iB�2ܨ�>���¹ ~�.�8�tFƭK��ܩ�Y�?̈~��Hu���P*xbߟ�S��P�g��^ȉ�A��r��_}�Ϲo�g�eq�ȑ��Vq]�����Z子��3�_���
�J�s���R�~6�����w���T��8�C�uv�\R���d:GT��-�����P�+���|:��ê\*����m��=���Z��-�)n�Ehr>C����.H�T�8������d1��xu����~ܝ�g���ȫ����YY�Ա0�'��ֻ8�mS��Үn6�!���d����e*�Ϸ�ÃM���v��P�.��KJ08e�h��/v��v�_��������8�dq��+7�	�����rs�1(YYt�7�b�v)�H�G{R�䕟$��%g�+=S�~s��s��9��%��������ֵ�ֿ[5q�W5q�Wԏޫ�j�ֿ[6�i~�iwy��K�Q�e��F/�#�w���5��!A�Q�m%��ԹO��x���1������c/AԮ|�s��#��a�k�k�ڙn˞��������V��fv�i�����n){K��Z�/ej����_S�K�=1Mnh��R�=�D1�q��>���z"u�X���P�a�/5����o��Q��Vh��G���s�d~v�?�v)����� �$d��}��A�J^�t���{I�����'K�N���/h��-��A�h>�K�Η��/[:��Rت[Kb�lU-���T�*��Rت[Kb�lU-���T�*��Rت[Kb�lU-���T�*��Rت[Kb�lU-���T�(>�٠�4f���}��A�h>�٠�4f���}��A�h>�٠�4f���}��A�j^�t�l�z����������i��"�)����6t[6+�g;Ԭ�G���u�޸��1������|1���Z�l�͛y�o6m�ͼٷ�6�f�l�͛y�o6m�ͼٷ�6�f�l�͛y�o6m�ͼٷ�6�f�l\m���q�S�mm���Ge>6ѵ�6�&ה��^Sk�myM�)�]��.������������C����mVu0:�
��/�Z�H9��H�Q)s��i$j~��{I����vU����X�H2-{�����w)(D�xd�|�)rJ��ku���Y�[��֤/��vG�՝mg�A���!Q��W�F�~Veߕ�b%`�e����:ȥ2P�l�6��is����8�:M�$�&��	�k��Q��w��+dTlxz쩝���|wY�y����Uh9Y|�JqzrJ��ku9Y	��і�����+��C��x�iz\��i��Ʋ�KSv��/:��\m���K�ܪ;̵��Sy�C)�'�h�lR?b���֥f�+5�SZ�5�SZ�5�Y�~��ef_��πޥmg��� �c�Ge�=���2Ge�3�g%�[�á�ܜ�X�݁��/F�3��z�BtBdnB�7.]�k,�L�g�r07,![��%�h�"��ۦ���ȩ5eU�w�K�U�Cx"A��qx1Q��-ќ�g\I,�Y�l7� ����*�S�ܽjY#��:+ �H���S��`�׍ͯ_cM�������R=o����.R�c��R=�"�<�=�!�~:�l�d�uJ;-�jv�V;-�q9H��n�l���>�o���U���ơ�%eK���a�1��x0�+��^�G�x��������%�l��?|,������� Ď���NC��r^��b�5����ʡfS����+��/2�W�9����)���,���nq���$.*n싕M��xWo�6;��\0����Ǣ��o��6��vO��iI}Df)#Ab���SQw�ĳ�K8�%f�+5;P�	Y�I�K��u��R?z��ԏޤ~�#��������������ط�6�f�6(cb�6/��l^�ݴ{���ŵ�]��e�{L4���nʇk/�m.�K덝��S��d��*�ML�\�1�W�yS��(�5��[)�|���k�����;|{;}kM/�������}o'Y��g|��:(|�q]g�f��/c������h����D�{	Q�c�r�ùO�J�E4ύ��#X���Y�S7h:�J�v^F�խz$���7i�����u7~5/vY#���b���:�ùK�)R�.|�KX��-b��A�S�� ���l�~T�6H?*%Ki:��R�N�A�7��j^��/[;�)s�.|��d��=���\�K�)s�.|��d��=���\�K�)s�.|��d��=���\�K�)s�.|��d��=���\�O���h��>6����h��>6���u-����Kb�m'Rت[IԶ*��u-����Kb�m'Rت[IԶ*��u-����Kb��n�䪴V8>��1������mmc�ˤw���^�j�������Q�kh���[ۿ���c[�g>6ѵ�7��b�l[͋y�o6-�żط��b�l[͋y�o6-�żظ�Gh�mm���q��6���6��ה���6���yM�*{^R��R��^�K�)z�/X���b������y�q�(v��O�vݴ�Hح��6��Y���Fi��i��s��1}Uke����6_u�]n_�m���e�ն���k$,�\�٥�FJZ�9-{R�y	�7s�eN�J���=2C�-�N#Q�m��yk�B�s{
�m���v"^B�Ccti�0v�ۖ�˿���R��>��VRT��[�B���*��Y>�=��e�_810�*?���-�bR�Iؾ�) �2y��E�O֧���l�6��}��n�{I�����[��F}�����W�661��J� �Nʗ��Q���e/L�e��c�Oԡ�3y�R��6���Oy���6S�6J�c<Wf�vl�b�v,�f��6s�R�/����;[w����kmd�k���H�8l���r�-G���Ӥ�M��P�F��x�~�9��U�Dл��l�4����p�$/:P\�9���&�drp��l�������@ܬ~`�%�?a���v�R��^�#��=�/l�5�
^+��xL�'a+=��2!Шʂ�`�*�ہ��蒲���7�����ж�j� Ǉ����s��������{���<���%�mK�����K��ê\/��Gm�x;��zX;�E%g�K���q�褬���U:�qn�R�4<VK�5�+%䵲=�ۭ�in=��k�?8�d��P=�i��%gKA���pb���_�J��##�m��H��e��u�^�8[�)��['���x�O�ò��ld+n.?@�¿ z����(��_5ƍ�W(_��G��UǶ'9��H�����VVl'+2��.��s�p�b��q�W�q�W�q�W5q�W7�g?����_��_l�\r��6S�m����q�S�l���Oݲ�e8>�R� �%Ke}/i���K���z�i����KS~�,�k'Ϊ9TeV)ʣ�.ygX��_dS-v���#l9�w�m���|��]5�v��S�J�\d������qlu15=D��݉�2V��H(�̷(_l�Z�e�e+�.�e����J�Պ寶k���T���>P�줫����b"k5�Mk)�Ǔ�I�o+�*�i��t�ny��t��"t�E�����⚙�5�~�pb��X��g �.z��ܥ�Y|;���/�r�=e��R�C�Hw)�!�)��H~�p���@5�� � �X�kb�@5�� � �X�kb�@5�� � �X�kb�@5�� � �X�kb�C�Hw)�!ܤ;��r��R�C�Hw)�!ܤ;��r��R��?d���!�)��H~�p����?d���"����ҭ�i=���ؿ[6+�b���f��=�ʻ�K�6|�;��{;�m�ƶ���v�{]�k�T�M�ŵط��b�l[]�y�mv-�ŵط�K���i~�b�m/��[^R�myH>ɵ� �&ה��^T����u�`���u�`���u�`����7Ե�^����K��R�)z��Z��z��=e��M��e�=e#e/��K�6tb�ؘ*�'��ʬ_(r3�	|N"A�G�ҔAJ�I�r�&'�aN�Q��z�s�2C�b��i��`n\y������*�%bE�Xȧe;r�1|��)��c��(�c��[��HZ��tw%���Aew.2��;8m&��ۯK49�y0�4$���Y�w{���V<�����*���������Ւ�X����jx��]�ž?#��fOK��æ�Z�d��1v|��Z2J���`G�=,@ܨ�Rj�"+��-�W�v��{IyoL��M2��o9Hce8cR��P|��2Ӄ�o��o��o���Oy�CK�[K�[K�~�#���I}�G��c��څ��<v����摲M�&��+dhso��ɬ73V�<?�ȇ�I:Op��w�8=���-f��Y�ѫ���3_�YO���J�W�����ʶ[<�O�-z5|yT���d���?Y�$l�����e���R�dujE��|ⵟ�vS���U�K ��rү�يwl`�h�V���Q�M�����ß_��b7d�j��<���K�?����W�L��Ge������S�{-m�R�j>Z��N� ��h>��OS��Ye/�7ݒ����v[�e�:�쇭��z�M/���61�GʻQ���������"�	����>����^KWǃP:X^G��9��lV�J�Vxd��/���d-*�w�9�B����ڣ,�[��U���%��fO�wd�.�����H?��V�^���F����Vի_�1�P�2�GnU�&O#�4����q�%�Wd����θ�_��X���{U�uo_�k��W7�b�l_��ط��i�e?w*�v�~�d����yH>�� ����S��.�u�`�����vYs�_s�U��Z��. �?�-o�R����ñ
�u��9)�K���m��?L�ΪX�{$��o��3Ht�L�˭�+v�("�k�,v�#��_/�[�J\��i��ԫ���͞�F[�y���U�J���q�"	�Fߝ���.~�m�LD��g�+��J�NF��9A��-v�N��Y�-�ˍ�[��I���e,�N�+֧�� �O��� ��tө�g�N)�E3��e�L��dS;8�Y�݇k/�jnõ�õ7a���ڛ��e���ٖE2����"��S8�� ��)�@53�kL��S8�� ��)�@53�kL��S8�� ��)�@53�kL��S8�� ��)�@53�kL��S8�� ��)�@53�kL��S8���_ �!����;Y|��k/�r��U�v�p�U�v�p�U�v�p�U�v�p�e�R���C�R���[�ʍKe}/i>6��ظ�b��U-���i|{iF����Q��/�m'K�N���/i:��t���[I��O���|l�}��d��%K���-b��T���)R�.|�ƥ�>5(~��C���J�\�vYs���\�e�<���d?L�gP�2�C��u�#�dSS|iF��߈e3���Ku*Eo�ʲ{�U�V�NB���6p�N�vH���%(k)��Y�Bod{<_�ݶ�E&Sxte5���޺lF��(b-ջ�0�o�T�_��vCc����nR�G��i
ON���$�_͌^2�������o�e��b:�x�RFˇ'%n����yW����t���R����Ab���lB����I�4��\��T�rZ�wYr�E�v9Xߗ*O�����u�?i(IV?����$A�Wƚ))o��qI*O��I��9��g�vK�j�=��?��-F߽��3�֤�w$�䥻$��%�i/��<���)z�{�vw<��Z��ܪ<nU^��6��Խܧ���r��*u��+;���K�t�&s�E56�8�=lV�Q�iV�D~�~
�����Co��}��1ޫv�8v���6�pRy<M��?(V�cn)�X����s���͟ggf��M��aY�6�D��vWrX>�d^��ݑ�L���H��G�b�n�2��4#�������I>+��U8������h�IB��$�*�4��?Q�����?9�<U-�@�Լ|��x<��:>���fq�G�?��+%�g���Xk��i{�1�q�����������%o��P<����$�B��rx>���0�՜q���+%�[Z�����ǀ�\��+3�����:�sn�{��9s�╬MvP��l���]g�����|<��������c�Pc��:��L	/Y��v�l���[۷�V�R������\�쥫��D){	V�Q'��i$�f�y��#����+��-{�,Wf�6���7�41�~���C&�d��}�ʞ�iwݱ�KΩx�����v�j[+�z�?S8vvp2睜;;8�US�!�*�T�OFG�咲HȥJmҕ��[�SM/S��2)�������HK|��e_i���nyj6�켷��#d����u�%�E�~���L�y�qy�r���=��R��6�l�eMj57�	#IH����P���w)���U��+��'wʔ1줫�}�kw����$i���-�m\\*�>����Yz�+��[��8��D�qQ�a��o��2+�Tq
�!C�(ze��<B��P�
���C�*y%NJPr�fuC�(8�L��T=2��P�ʎuC�*9ճ:���ꃖ[3�YlΨ9e�:���ꃖ[3�YlΨ9e�:���ꃖ[3�YlΨ9d{-:��N��G�ӡ�Q��z�{-:��N��G�ӡ�Q��z�{-:��N��G�ӡ�Q��z�{-:��N��G�ӡ�Q��z�SS}�Y8���f�p�U�*�?�v���*'���|l����C�S�l��N)��Se8~�p���8~��ʜ?d��N�|r��>9S�����O�T��)��(����C�3�k�L��?S8����C�3�k�L���4��� �#�dL�i�2=�@4��� �#�dL�i�2ٝHx���Eu*��^+��O�F�2������OSvݦ���Uru�� �SU�EYm ���%׻[ǲ����j�w�d����p��ek�����C�\�e	3{[�������ܡ�m��q[d�YVJ�~Y}��"~�m�5�$�u�o�Dɲ��"�m}�B/'B4V$���>V�R�,���)�Y���}�pZW���%�U�6�@��v[��=�۹Y�H1[�Ǖ���_�Ʀǳ�p�%���=go�%k0r��+����_%?D���Z#�8���{l���vxq2�H��oG�^�5�;/ �N���Z����KSw�-}/S}/SR�k'��=���6Ov�\mv���o��I{�[F�SX�J�m�OeA�V�4���Aה?*���c�gU��:<�}�Wj��i6�Rl�U�A���}���<,6�2�>8*M��ny�ڻmܯ�kk��^�e�P{�0z�V�#B�Ys���J��g���`�V�"��N��-��~V�K�i�����8��+����%\�9Wz�� �yYmNRm�D"��ݗ���۶�f_'�Vb�4�s����f�������֭Ժպ�Z�R�;!����;��W�R�[�u�=+(qIZ�R�����[�Hu�b�J����L� �־(p�:�s�.;�V[��>�K�[�����|yY��62�)n�>U�D7���������n|z,���/L����J�/�n���z[=5;��W�t��O��[V��ռ���)�Y�?��� i{<��>�R�7�:�^Sy�b��h��8�D1�~���d�r�mc�X��N��;���gsΩy��eV��S8�Y����)��)���_C��<���l�ڮ�p�5|VFώ��S,��ҕ���/Ūx�NJ�[�Վ��u9�9l1L�X"q�)S��L��zm�*�-�ݦ���']�F[+8\�_a���������M����J���n}�Jyy	L��4}A���b��6筐c>\�TC����g�V8�X��gZ�\K{HH����R����%��	��F��C{���H9�R�:�����ߝKzd��Etʎ!C�*8�+}G��o��<��B=��Sʪr���Pd��q
V��USʪx�O*��<���T�!Q�*:eG��B��Tq
��Q�*:eG��B��Tq
��Q�*:eG��B��Tq
��C��C�N������;}-:v�Zt4�9�M:uA�N��PtӠ�T<��<��y��yi����ӡ�o��C��C�N������;}-:v�Zv�M��M��M��M�R�@9H) � �������;��r�=b�\����s�!ܤ��k/�r��e�R���@53�kL��S8�� ��)��S,�e�L���dS;8�Y��=�E3��e�L���dS;8�Y��=�����̪��[2�!lʨx��*��̪��[2�!lʢ�e+:��J~!Q���#m��ϖw��B����n��Q�U��0֩��)����Yn.ԅ��ICF�A�ʈ61���Fߕ����&Z�ַ����u�"��o�	��h��rCla[od��g�a�2^'~Ϸg!K"���69�9rl��-g ���I�;�X���d��A�5�J��=Oeʵe����~M��&�o�sȄקg�P#ls�,�V"���iS��!���
O$G����/X�G�rv3-�������6[t�~.?qʠ_Z���rUd�~S/���:nz���w'aL�R[�v
՜[�����U��S�eo�b'�_�����Z����|��z��z�S~ה��>2��Y��o��7=d'++�(I��z�O;�Sk��p�ִ_&�Fu�������QK�]�V���ů1?{5t��D���p�I�u8��:>���$��80]d�Q)[60��KJ ��-�-�������v�_c�s�`�xi m9�H�h��q�ߨ��ͭ>S��~ݞ���?vE�)P"�������Q�Ⓑ9�emq��i#�8����!g������xY��0�_K�x2;��g����d��9����<�ޜS���,��으B�qOS㎡ó���xj��qO��=��+n{Z���tr_8�R�?�%�l�� ��W0Ď��_��K����Dz]�����6v�l"�
^�_#K�g�
��2!���Z�H�o�>�Ys�v�+x;<��V�:��Us'�F�|���<��E]�mý��lNEK�c��b�5����C�-�6�F�{��o6O���h���S��o5�6�R�#�dY|Sev��T�{L�jn�e���TB��G���4�c�j6̭�V���;|���mEs���)xwv����b�e1z2��2J^���S���*4����;qL���Y*2���
����S��R�9*�/-�C��y,�쭭��L�s��e��˕���ܔ>\[Mn.��B�<FmD���n���rٖ�$H^rW+�Ztf�����!����C��iR�Oc����$)y���ݑP~R����i(h��������F�$6�^�FC�N;�V���!��)�-�R+���JErS��H�Jv�)Q�ݷ�J줖�J��|W}NJ�[�+�Y�q
�Vu�B���w��g]�+�Y�q
�Vu�B���w��g]�+�Y�q
�Vu�B���w��g]�+�Y�q
�Vu�B���w��g]�"���dW|WL��/��\E�]2+��+�Eq�tȮ"����_�*zk�<��zk�<��zk�<��zk�<��zk�<��zk�<��zk�<��zk�<��9k�9k�9k�9k휥��k�b٬��Y;f��f��������Z�~Z����2Ӄ��S8����������������������Zq���iǲӏe��N=��{-;fulέ�i�3�f�v��٦��:��=2��P��!C�(x���T���Pr�UAʨ9U*��T���Pr�UAʨ9Uw��1�4�d��e�J�h��Y�R���jʷ�
�IQ�ݭS[>��emWu��h���Y)h�b��+��jrU���V�!U��6\�Q��,e	�����q;�lC^֖���ҁ�2�L~��'��ӵ�Ф���Dݶ��)��]M�M�,�یݔ5b؇'vX�$�n�+���l�y"��Y�,)�h�+�l���R;s���N�b07���S)�k�n[S�%z!Q��_�c�ߍj�e�;a+z��Q�d�6q{����w%FC�s����{JOl��e!a��u���ζ&+�����4����9AQ�-�[�[��R��L��gs���-|-8>Zp|����2ʖ!�� ��ԭ�Nw{��B��n-���nT����q_�����Eg}��0�K޻v�����rh���:����[-՘1���9c��P2�=���;8I;��9!�y4�݋��؉*F�۲���/w*Υ���P,�Bu�֊�����4��*��x�?o�Ü%�WvOg��*ȍ��AF�v?,��jU,R�l�h0��絨�5@��1KuO�����?��l�[����1��@6��j߼�)[^�^���E}�8�R;�־6>��WSL���LF�H�kd=��[��j{݅G�����#;����QZ̑��{Z�G����9�A�e�#���VGJ�_��9oiM�R�-��*Uj�U3[�S!T=�|1������c��ϖK_岦�?;-c붋J��q�Ѱ�Ca��J��ۥ��n}�v^O��ld���������b�:K���Ke}�i|?e:��Ը�f�:�gP�L�x�WS:�*���S�O;8~�ճ*��TB��[1m�Z59*��|�(-��T�}�/n�K�$)z�
�����q�t�d��9J�A�@����K?M��{l����e5n�����=��񴉊J\�nw�H���V��
_/(�ge�-5��[� ��s��T�Xl��~W4�NV�ȮJu�]�"AÓ��$mfEk'��)�z}�c���� m�v�AK{O4>Wܥn�w+�C��i�����+M��r��j��F����)$��H�-�%vRT�$�)%�I-�InRKr�[��ܤ��%vJ�[�����%vJ�+��o�NC�ܤ�d�ܤ�d�ܤ�d�ܤ�d����9)o�NC�����9)o�NC�����9)o�NC�����9)o�NC�����9)o�NC�����9)o�NC��ܬ弬�Y�yY�r����g-�g]��[�λ�����w+9o+:�Vuܬ⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋⸋�zk�<��y�����b��T�*��S�*y�O:��V�4�؉Ǳ�en��a�[�D�i�tӠ�A�N���M:�t4�8�G��B��Tq
�!Q�*yUO*��S��U9*u<��%N��ErH����Y)�"�R+�ErH�I�"�$W$��\�+�ErJ줮�J줮�J줮�J줖�J�+wSFC�-�RF��zt���*���InAR�+�2�#-���W\�ܽb_%N���������xh9,�9
�Ki�[�c�C]�7��;�K;*�����u�*�I��ɤ���|P�鲭��l����J���*@�n>Ӡtoگ�Rp�\��C��J���o8���TbY?�y5�_~鸨�6~u���>t�%W)?���]�Vܯ[/M�G��������Cn=��t�L��!�1��J����=�X����M�Ks7g8c��t��u>����1��U\MaZ�Ѧ[e�X��~vƳ(y��П)�(a�So���d���Io��IQ�*9%FR[2�fU �N�@4˞vw<��Zi�ivZ�KSv�����K䵞nZ�\�A���h塪����j�l�ʒ��/���Y=[Lxp՜�5��X�s`�����9��}..-/1?k�X8b诂K�,9��ܭ?)ʅb"9jb)��\�����\��t�������Q�۠�b�9/�����M��7�WW�Oa�_Ig�Ma��l�t=�j;s�e!ڊ�H���ڞ+�b�C���ئq��?wG�9{�����q�����˟���?>��p>zVqު�G{!������,�����_������<����?V�j/�d�s��� �^I��"�>�B�6Z�}<[��~��mx�A�|zٰ��R4�۳��X�uQy�d��v�򙝓û�q�U%w;c�k��<8��@�ۣ/.Nw˒�p�%�����zn_��� )/Z�@661�d�+F=�����(�wbqZfG-��ʫ�KùWa����ʖURʡ���4ӷ�/�eR���/Y���E���%:�!Q�*9[�rU�YJ�9AS�v.��.��W)!Q��j��X�JaX��D�2WD���������jfZ6ى׭l�$���앎;!N� �R�)Q��ԩK���/�� v�]�KFJ��+[�!�3���܊�[��l�V'_% ��b��d�r�bt�rC�Rܥj�)\S�2h�'�H��6~؄_F.B��J����P�{���aQ����"�IJW~�qN�b���/E?��e�Vʎ��F-O��ũX�*PR�h�-ţ��w����Z;�R�+�҄�҄�<��~V��%Q�JW��%�P�vR[�	�e%�P�vR[�	�e%*R�ݒR�+��%*R�ݒR�+��%*R�ݒR�+��%*R�ݒR�+��%*R�ݒR�+��%*R�ݒR�+��%*R[�JT��d��In�)R�ݒHy)Ҥ��y)Ҥ��y)Ҥ��y)�y)�rU�ܕ|�%_-�W�rU�ܕ|�%_-�W�rU�ܕ|�%_-�W�rU�ܕ|�%_-�g-�g-�g-�g-�g-�ޙ-��2��Wq
�!]�*yUO*��S��S�䯠䯠䯠䯩�S��S��S��S��S��S��S��S��S��S��S��S��S��S��S��S��\�+�ErH�I�"�$W$��J줮�J줮�J줮�J줮�J줮�J줮�J줮�J줷�|���|���|���	PGe	��{)yo+:d���4���:��M[�e5Z����M4)��I��u;�N�����U����R�$[Pl����(r62���V���ߔ+iI([lk�����Ȝߔ��,:�p+�fE�Od~;N����۫'�X�V4�{p!V��C����eR�r1��أ]a�8��N�j�}�m�����4e��eMX�m�d��ևʇd�+X�>�m�������jw76qyf/n�E�!kӻ��nG�i�������Xַ�4���d��H�p�rP]F�C�`e�z��_��v���!�b�T��R�-���-]��\��r�+((rR�%#�R)�E1��>2���Ux�l5-����_-vB����%[�y]tB�_��n���@�m$��.����7�$�j��ݫF�5�����6&&YIa٥���������r�Y�����K �W+8-ZM��a��b���B/����G{����Y��l���J������$�.�ͯ'�����e2I��	#i����ғ���.�Wf;��A�v�)*��☤���c��ҏ��YϏ�ǾK�ެR�t$ܩ~�o����^�$w�8�;�ǁޮ3�|1#�����b���G{*^�b�.�K�"�.�K�*0�S�i��վ�+(0���j0��~)},y�� �}>�#�58b�]�V��?��H�l%�ԗ�a|��:���b�%Rj���4˒��݆�����D�����*<�UG{�蒹=�IC����������
7�3l��j�K��R�X7�~K�Y���j#b�lu��)*�d��yڶ͖;g*�SM|zJC�$RRP�W�r�e��]D��r�[�_r��ṰYo-����Q�Ѩ�o��o��[�Ε!N�!N;!N�(]�d��R�M6�^�WQMѓ�|�kz6ƢB�#HY�k.=En_�M͓�Xҽ�����H�X�q5�
�>��V�D���n�u0Y=M��Y_
���HZ8���a��T��o��dT��RR�{s���l]X����e��@�+��`m��
��_۝�����,��*�=l��Q%c��I�����M�-�S4�4��;�[o�Z�Q�)YtS�m�U�ʧ�U�,��۶�v�*�!)��!)��!)��!)��!#��w�J��Wm�Z�ܕF;�I
��S�j~-Oũ��?����Z;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;(N;)#��;)#��;)#��;)-�%�$�d��ݒ[�KvIn�)R��))R��))R��))R��))R��))R��))R��))R��)$<��9)!�IJ[�+�����)�rS��\�+�Ed��*��V�)!�JVUJʣ�T�RT�<���)��S��o�Nߒ��%;~Jv����)��S��o�Nߒ��%;~Jr����($9A!�	PHr�C�����($9A!�	PHr�C�����($9A!�	PHr�C��Z��R�jV-JũX�+�HKu���k-R�����-�[�����삎��9AO����z��/��caN����c��B�-Xm8R4^��e����H���F#�o������c5�mXo$$~�m��E�q��n϶���������kI����r�*HKl��"������Q�Qe�y))#vG�D	ic��Y�~�����$�ly���Fj�Yܥ��	�v2!���4��o� ��S����A���z�!(y�# �cr��*����ZRZ�Yݷ�u�6+c����6�~.6ʻ���S��wd�j�����W�y+�ܡ}*BR�%vRErS��Io����%(rR��[1�!ʢ�U�d�v���� �_!�T}�XnvE
����j>Y-6ʛ�Ҡga�݆"�L��ܬj�U����5�pո��M_,�B��>Gp``k���Z�O�H�L١�Rm�Z�m��y)�R��
:%�g,�@����)R��p��V]o�[����BASv�����(�d�L��3��D�w7YI�����Vm��N���2^���8���Y�e䊕j�\V��Ƣ��Td�j�\R�9�F�T����%������H���ϏEf!��dR��Pn~=F�[*]-N��`F�T���=�T��P"�.���~$���h��K����-�y[*��G������e��X��'�݇w{��b�}���܎崢���϶P�`i�q�-��5q�:����;�ݵW7۲����W>�e�J����<E��K�����
~"�k- ��ryYz�ǭi����l�]���	C�J�+V��ʹ��<��"EO����Ud�6:|�V[����Kt���Q�!�WjrU���E�+jߦ����l�q5�Yz�m�o��A�_�q�$��4���N����i�1;,nJ'{(y��X�4۵�j�eV���#�wg"�G{t����L�f�'*E�]�����6�$B�M�v��n���zd���m���V�������ʑle*L�6�'��j$98�ܜ)#D�ڵ)12���[aMe��I})Kn籁�`�e/��-T��YU�j;[�[�]��w�d�eIT� ��$H)"AI
H�RD��YU�*�!N�)Q��y%V�!O)[V��ՕZ��VUjʭYU�*�eS�)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��jԄ�HJԄ�HJԄ�HJԄ�HH�8�8�8�8�8�8�8�:T�}*R��)_J���JWҥ+�R���J�T�}*R��)_J���JWҥ+�R���IJ���IJ���Io�*��*6�J��R�o����S��o���)!�JVUJʣ�T�RT�Y֤�Ҥ��y)��+�Jv�J쇒��R�!�-�ҥ$�(_J��ܡ}*RKr��ܡ|������������������������*BR�%*BR�%*BR�%*BGqh�8�99;|���|���
V-JũX�+����Z��Gd)�2Y�Z�J��/e鳮�lm��O�~��n�F.��%�/���Wc�\���^C�ڷH,�-��g��e���|�2Q��n���M��c���P����e�_�%g�lu�nB�I/����^�P�./RRuW�\B�V��?z�Q�ҌϹ`�V9(�o����F�lq�4�[p����c�#���l%�|~��fD%��������J���Y��~�/a�@����r2�'�$_i�!��m�Ci�ێ�t	#)���ɶh�L^�c!s�B����+kc����K���26"�2J�L��O���HWm�[|�F[�/��jIA�-���)(rT�9UL��5YP[��k'��a�k! �5OY���ȤnUb�m׉��Õ�b�RB�r��Ѣ�����MV�[R�y�D����5��5$n�:>��&3	[�K6y_��<q�-�فg������O�f�+[�ʶ4��N�
���@�\Q�U?Fw;+x�Y(J���)>�ՓAp���vI�c!+���Dv�K����?wG�x6ʗK�r��@�x�
�Ik$��z|��>���Y<5�q��⿻����3�|��z|i/ԿR����?�+��\g���|~�Q��9G8�;�Ď�|C����><8�k��i�c�d�)��\q�:��$e"�-EG/$E5��"C��8�Ԭ�V��9|�_,���{k_*���&��u�X��'+Ź����&��K�WŬ�ڝ_�<D6#H2ަΕ��J��e�"���x��;�Z�k�!a�H���%.H���.(:�TE����U9
uB�w%V+ʸ�Gڍf���ٔ�Xr����k��W5jP��ee+j�aL�Ο)c��a%��M+;q�y��2x��9����y���+��e��i�)��M���+��I�:�������kkx�T�8���enu�,�2B�e�5]6��@�T���^�m�m%U�
��k0p52(���P�=��;�{m��Z���=�-���J���S|�-�2FvO�Q�[n�qum�*��+�l��D�/#Yn�aO�o]�V�񱯒�yRW�ԃvH�T�j�[I���e:�e5$SRE5L��i#H*e5$V��jF��2
� ����J��%a�d��VY���2�:e�t�,�VY֬��YgZ�εeV���YU�,�VUjʭYU�*�eS,��YgZ�Ο εe�j�:e�t�,�VY֬��YT�	L���	Z��R�!+R�!+VUjʭYU�*�eGqw�qw�qw�qw�qwۥ	ۥ	ۥ	�e	�e	�qw�e	�qw�e	�qw�e	�qw�e	�qw�e	�qw�e	�qw�e	ۥ+��%�$�d��]��Bv�Bv�Bv�Bv�Bv�Bv�An��I���I�'Z�'Z�'Z�'Oũ��vB�?��S����
t�Z;!N��Gd)��h�:~-����O���U>ʧ�T�*�eS�}�O���U>ʧ�T�*�eS�Ֆu�]��]��-�ݖu�	����!-򂕋[��Օ$H*e�u�]��
�v9?v����)��IX��[e�����uk6�nʃe�Cce	5'l���_L���Z�k' ���~�v��ݬ���Vv�[�qd�"�~\P!�{tҬ�s#dPvW�m���Y�Ȥ�o>�4��Ќ�is�d7!3YeR�Ě��ڽl��g� Z"���T�iT��Xi���_tj��ȉ�'�F���E%ń$n}�}�Om�v�}���F�{��@�{Q��wx��#-\��rW�nDȸl+y��6�Em���JP��:�Q��҅%6��'ݹku�;M������Н�L�H�0i��Jַ��MV[�FGq98l���U���;��!#�T:�;d�8�.t�In����[�a����xu�9)�Z����T�)+#Kw�;r�R�o��K)-s�v����e��E|�Ύ��汯����_a&�Օpܸ���f��{��rȸ�D��@Ҳ����R���Sk��KM�Z��ǵ2xc'�!m�����k�f#M#l2��<
J�4dm���*�����ξ�s_������pb�C�n{^?�#�Ԭ�~�g�K�������^K{!���|	[�|�+�{���g>�/�w1HY���q��󎗧�A�_�w�\��Ƒ��/�+}?>���W8��;����|o��������cל���9�q�w�9�>;��J�:��J��u�;��[q{*m�;���h�);��.����=�]�;i
��8����k{!{d��c[�}��[\��N;�n�E�r���x�18��;���%j=%K��<�~';��Nkl�b�|[���*2Jrܡ}vP����S����S��S��QܕF"_����Z�L�����J���B�Z�/�IX�]��7Ev�������°����e�wY��ףZ��Y.IykSN�]����;.VZ�o[I����d��+����學�0�Q�J��F���t6Pû��[k�V�ƛ�V'S��������o�T9M�
�- 㐷�*����;��R��;
�&���[����~VXOmoF&��'m�mH�En��^z���O~�ӷ6A��jpc��=b��Ye$�e[�	ۤ��,yNW݌�/�+���v��V�
kaMS)��aY�O/N�v�w�N�Y�O)X�f���՚r�NVd�2����6��6��6�"�|� �����H��H����2��SR55���'M��[�>�9"�|�[�'M�N�:ent���jj�ebl��-Z���	$YRD��$� ��) �������ԃv�e�>A�>A��ʷYT�*�eS$%2�:d��YgL���,�) ��VRAe,����YYI������)($lZ��S�j~-Oũ��?����Z��S�j~-Oũ��?����Z�eV��ՕZ��VUjʭYU�*�eV��ՕZ��VUjʭYU�*� Ο Ο Ο Ο Ο Ο Ο Ο Ο Ο Ο Ο Ο Ο Ι ���h��5��A��A[�ʷHH�-Z���*� �T�R�~NA���p��+�/G/!@ӷ�ܴ�C�䲲U�n��ɤ)Y����ժ�$�,��Ȣn-��z���6W����;+aNobl���թ�����,�7�vB��Cz��q=�iU�������r�,C��뿻�^YIۃF6�˞�m��$JI~�k�.pZ��cs]��GWퟢ>���h�cd���mOg��U��Wl4K;eZ��)x�ԝ����~�N�7���J���/�����y�Ƶ���ҫn�/��G�]�ܽ���l�v��L��	�e�;|����S%�Ke����ߒ��Y�m��
V!�E:�n#7+W;!Oc[���R�=g�C�W�i��l�nBTl�6���}�B�n�'n���)��+VUG+|;;?��ʣ���vq�G�JR��xd.��Tnޓ�?��e\�'/V�2�pᾍ���ѵ��#�E,��XBW�Xʥ��>�B����Th���K�W�$�OO�}�Yw6Tؽ7/����~����ۗ�LٳQǚՍ���!J�Fw���/Żß"�qJ�$�:�#'n�`������^������OϢ�{�|��C2[��~}/���,{�~7s�{���o�� ?~���o�� _>�B���)[���od3\��l����-���������x�q���g��<�A�_=po�-��R�K��x1��y\�ez�ҲV�)|wgZ�l)T��o����6ˬߦ�V��P��+c��j5��O$�e��o���0y,�5���(Y^��«��USM�7�&������9�,�1�+ͳV�)U�� e���^J����50�͜���ק�Wm�%*R��(N݋��!_�ΣeC��Q�
y��J������#^����i�k�;
�#�����	}�;_c��v��^��\���'����D�zl�U˞S%g�����$o�$�(`IR��d)>�c��ݍ�G�ktNJ��jd�X�=��&���I�}D)��h�G����J�el$kom�B�l�i$�?+k��\�����f�J��4ژ�B��)���_+@��nK�)�Q�d�/���p�e@����Co��[�m�o�ۏ�����W��J��iB��� {����/e-��)������d�Wc�����9L�>T�ʚ�V'��)X���]�Ө�i�k5��J�ܽ:�^�<M:x�t�����u��u��j��5n�ent��镹�+s�V�L�ΙMH�ԍMd��V����)�����)�djuEn�En��:t�u�5nz�����	Z���U2��ST�jF��j��j��j��:��Jmܥ6�M�H��Z��T�vAV�2�9�9�9�9�9�9�9�:̂��*̂��*̂��*̂��R6-�ű2Q!)��!)��!)��!)��!)��!)��!)��!)��!+VY֬��YgZ�εe�j�:Ֆu�,�VY֬��YgZ�εe�j�:Ֆu�,�$H)"AI
H�RD��$� ��$H)"AI
H�RD��$R�~N�~N�}2�|�[��[S)�Aj,�����R4��+j}:t�u���e:��Y��Q�e�t�*���m��Gv�"��_/�����
Ϸ�n}��:³����Z����i��m#HJf.�v��γM���F�v;{
݆�!�����1�Q?��־��E�6Z���l�6��c×�i!�x(H�M�<2W�"`ڄ���"1��f䯹Gq�-Y�d���E��e���'��}��qgqa�c�(vY�6z�,̖o':O�M,��%���'�����d鸽6�l7�#����Jr[����R��+6��L��w"B�����{l^ԅÖ���H\���<�+5���H\��܍F�s���m �ػ���2B[�Ҭ��l�Ҥ%NPT�� ����<�����TSMF����r�$m�^B�զ���-��Zm�T���}�qڣ��\8o�E9�;�ݫj_���|��u�����&�g�܈����D6�93�ܤ�Y�Ƥ֬kw-�.�o���M'��)"��*��N�|lm���d���!z6;<�4��#"�rݏ��Cv�p,#h��.K�}��>}/��<��?<W8��ǾVqެ���/O��_�V��g�K���B�i\��_�#�Ԭ�\���Hu/Z���v���8
����J�����-�l�j���9��3����T�ZUF��T�T�k#[���[���UG���A�;~�c$z$j����r���w_���VUe��}��W�A�p#��V�PՏ���pȾʩ2��G�vJ��w���l8�9�FI���D��u�C|�+򕋴*�G%/S��������h;;��
���Z�/�J�J֥��D�|v�}�ʩ�R��k-@JR�/l�g��I,NS����V�6�2B[���؈݆�EN�V����6N�q����8�l\�)Xb+1����F�k��9.ۉ+M'�V�2U�l~_i!}��p4�Y6�c�L�ʶ0��b��7���6�W+�����&�o^; �T�(M4�K�����J23���r���oĕN���9nV�.?���VR�é�\|�/��u�D��'!h��h��yR]���P��B��5�!?�:��c�헬D%�1y�a�ڥV��>��c�W��WQ
I�N���ފrH���{�{����Ebw'�����_��_�_�_�_�_��_��_��5�N����t�4��i��9Y�15�&����zt�4��+�V'Y�]��.�)�v븚t�4��klMm��R4��ST�jH��jjF��'M�N�<�6y:�����:��:��:l�j���2��)�e5��U�Y�U�Y�U�Y�U����t�N���Y:k'Md鬜���j�-�ű2�)ee,�������VR��YYK+)ee,�������VR��YYK*�MS)�e5L����2��ST�j�MS)�e5L����2��ST�j�MS)�ent�j�[�2��V�L�����)�ent�j�[�2��V�#V牧N�X���N�X�2��V�zkaMz+ommY�2��2�:ն�R/wQ�#b<�5��v����2'nK��)D:�ړ�Fn�0l�?�0n�1��m'����jF���kk4۲D��)��ʅ2�7rr����G/ �i�0�W*��9n헒�%�}o=ai�cq)D?Үv���
m��&���@���.$T���W[����T�r��f��\Z�j��3�rX�
��F':L��;)���m�m��:������W4l]"�I�J����B�ȷ�i�ھ�X�:/m���h^G�2ڈ���r��޳_�Z��i�ݖVE��󔡸�VX�*�����od�-F�7M_�
�N�I��'��I�����7���T��R�u�C���T+�=%c��g-��
v�
�>Pє���r��B�c/�rE���ݕI�f�wtf��\8o�E}��to���+ߴ���+	>��L�ǭ���E;�-m�jk��#o��K�in�G�T(�$^R���V���V)��[���V��]��	5�_���+��g��ȕQ0e��n"z脸�a!H9)��S��N�$T���v�/l��h?,�QL���-E3�$T��9YA�p1�YS�g�n���yKw;]�12EK/���v=N�[�ld=n��A��L�o=�������yKw�S�b��R�S�c�Xb�S�Gb��j߼�TUt����VWb��K��C��v�H�巴̈́�A�r��,�7p!��]-�@�Ȳ~�n�i�%H:^ܾW�A�V���N�%�V��9ݣW66���O'�X�Re��.Fӵ]�\Ky*�ܮe5���9+5GS�[��ҲY��\�\���VY��Y��)�d�
F���Z9|\��B�)e`d�l�;����u��<�a#V��*��R���!Bi����h�6��BT���]��i[�[���m0i�T�F�p��T	B!��/![�[v[c�Ҧ¹�yZ��P����Տ�� ���O$6�'�FH�P��?*�i���'�?9�Q�{�*O�_!F��6^*dC�)��k�C~·�%(T�?�eі�_��_���ӭJ\.���#�n�>�n�
A�����G�b�Eo�?<�n�� ڥE�ۨ�9B
�ʓ��P���^��ӝ�l�yۡ��Co����G���o��������g��OcX���=�}菾Q��>�E��Qj#�a��5��S�
saN{iͅa��2��R��[o��/�ӯ�V/��Z��QXj)�Mm���U��Ne+lMm���5�&����zt�������ӧ���5�&���՚j�[d鬝5���'Md���Y:l�t�N�<�5���'Md���Y:l�t�RʦHIBd�&N���Y:k'Md鬝5���t�N���Y:k'Md鬝5���t�f��ӕ�r�NVi��9Y�+4�f��ӕ�r�NVi��9Y�+4�f��ӕ�t�4�f�:�9Y�N�NViӬӕ�t�4�f�:�9Y�N�N�^?<�~u��F����mVm��a菶�&?<���D~�/w{�e�vB�N�j{��v�6D�܉��ʢn]�;���V}����6��X��\����v�~��G�(s���l�*�����%~\k#�a�
oc�X�)~Z�� e
ĳ?r��GrOa���V��[��'r��=����9<�"�|�+�&c
p�Q���phO��O��éյ)g�֘٫��g����oӵ䭌7+��v�k��a �97)��{?8�0�P�xi0e	C�ű��jv�n����v���Vv�����0m��0�,F�&�����[-6�&�����r�*�FA��966ߢ;�e�9��p^�~�O�"�V(֭�i��2E:�"�}j���QZjC�%�����[���n����NB���s�m��/b6�M9T������G����ݫVwn��to��F�}y���v����/�_����H7r&23�;��.u�ĪA��56]y~Y���wm�1N�E+ec����t�I�Q��})6�[��c��|�OI&���n���,wt��dX�N�8�8�^��x��������^�Q�:^�)<<t���Gx�s���HY��J���!z�G{6�Ė�A����é~�󎗧P9x���O���>{���1%�����}s��$��Vx�R��K�J��B�/G(�^9���>�#P%l��x=��xZQ������@�޹��俏�/�x���k������.�D�r��C� �V%�-6�.P�rB�i�h�����e�R)eڵa.:�M2^�5�Yqe�Y�?�8�۽�.<���/MT�7�TvJ�o�c�b��T�6�J�j�:}�!�3�V��So�Sg��ߨ��[�,4�*�[ ڲӰ�e(/�B�GY{aJԂ��YHS'���\|����o���P�gm���ņ';���a��~dnF��@�IR�*�_��qS�	5���Ǿ[�潯n� ��2ػ:�]dC�P�!�p�[�Ɇ�+��K��em?����9M�j���-���c�Ó��O�Y���{�#�����.����/��Q����\�;7$��p�B�Ͼvi�ڵ�����H]��6V7��P/����P*�!R���đ)D쬰4��v��[(�[H�>������[�����ػelb�l]݆��ע�Eވ��{a�l5����m{m��a�;��v����l�1��c����ϻm�Ʊ=mb~��ae����^�k'XS�}���6�°�V
��N{i�m9�=�綜�S�
�a[l+m�m�����^�<�m��O/[e�����zt���^�<�m��O/[e���ӧ#[o�[h�)��5o&���ؚ�[bklMm���5�&���ؚ�[bklMm���5�N���:�'Xd��a��2u�N���:�'Xd��a��2u�&���X�kmbm�M����6�&���X�kmbm�M�����׶�?m�x�jF��h�F��1�&�����/@e��}�{��ܴBzhSem�m�Sd/2�Z�����,$(�(��e�`����K��~�vw{N����+��v����rU;�~�d�nVE���"���e �b-�u6Y>�r��xi4B~dj�d��s�@��rX2�}ĉ�@�"�O�b7v'�|e�n�~�g��h�x��|��`�ݗ��nխ���}�դ�oʾ�F�iD�%�Ʊ)m!Q���'��{7,��k��?����rg�7r�U�������ȷ��<�qZ���{M~�'����7>c�ΎEbE��[u�l�%iYd�VW�È�V��BP��p�11��ܓV�0#�1�B&P���E���5��e��&�<�5O��:�H�%�u�U:�+�k賖�ԛ�����Z�k9+{�dP�_�JO�k�`�%R��e��k��_|��v^��n΍�9��yT��|O�n���[
U2���qi���@ݍњ
ԚY�e(nHڞm��M��X���`��TwYc���\��l�c98xqm������wwr-���U�f��m�^p�Y-��p�u@��*�㽛�\��:�C��8�q ���K���$tV=�C�~v�#��9Y!�d�v�\V��b�o�Hu/]�H�N��]�H�n�����N)�Hu/���=��t����=�v+���#������G�tn����?վ�%�0�R�l�d�ok��ë6뜇l�@8�?��R�{͗�;[�m>�K4���[�!p�%��
�!N�����"?��q݌�"T4U����漼��ύ�rR\�/��Q1ߖ�*�GgN�����e����M+q$S��G�K-Ẑ�$�N��X��N�/N�ݭ�����"�Mb�&��g[��ea7�)Ki&��|�x��[��Xe#��+z5��nJE�����d�t���فGMe�S�9[<�v!(|��xn7dJ��\�*�{��
�M�܋ܡ+?*u3/ �.\쿗�*�- ��Ch��9�rteK�'��5�mn�*�o���!�u�0�-��v���E7�e,�+�����'��Y^6��/���J�ɶ����UVV3��\�q9X��JY,��$˸7tg��Ţ2	�M���y�<3��o�~]��tl��=�{�V�]�D���_��50�*��HS
|��ʠ;�v���[Hk{wh���;�v����k�|�D]苻�wv>����ckc�D]톱0�^����el���]苾Q��>���+l�1��c���g���m�ʰ�V*��X|��a�>U�ʰ�S�*s�N|��a��׶���^�k�m{m��a��6�°�V
�aX{m�v�z;(�=�o����aXl)ͅa��6��V
saXl)ͅa��6��V
�/me�~y{k/�^���痶�����~y{k/�^���痏�al"�]���v�.�E��al"�]���v�.�E���X|������1��c������c�����G�@���]�v�,G#���]��M��?�%`exn-�.����W[ѓ�\j?.�"vu�rTB�-�%D(�T
5�Zmc�6!ϓ�^�����`Y0�y.����b��\�����I�2#k{�[t�;�w���C���^��ߑQׯ�,�����M*��ȓa���cf�w? v�����S����%~m)[\6�,3��	�"��ҭ���{dR���/*�Y��RyȤ�Ń٦��>Q�V�^/������v���W{v؟n��m���26�[���K#���&K�A�G�8��wv˰��Q�^�w��:&Ym���_��o��<�9,U:
��k[@ǉ�K��z98�݅n*k[e)�u6�w��M�]�AR���M�ʱI��m��MO%;n���ݽ��m1�V)��c�����ݫj^��e��j�d�66Mc'ҳ�9RVN�$gv�lB/��B����%XȈk��Ae��rޢ�!v\m6�+���*�a�J��i=���!vF�I�7�y2y:��i�����K"r0l<�Z�����'����~QZ��o�l2�Ol����;/E�e݊��p�����*[?m哀Gk��j[�2��5f�K���Ze+y$H~�;���,L�R��$u����t�o�Kt�l��謏�|B˟��b������ø�R�R�K�)�[K�J�_�V���#�gώ�z���^z�pc��W<�A���V�������#e����ܲ�x�����rR��vE���g�Z���"ȕ^U*�:7�&��U�*�fܕK�s��}g�g����2z&U��+�(B͔���[g���H3�SgO�_�ݦG��-�vv�;J��]��߱���G��5�T+g��n=���k'��=�{�{/�M6/���J]�؅�ʳ���l��(/nN�)d��nVN�����M⸋�c��k��˒/,��[zjn�OgN�I[u�Ȝ���[����>d[�o�J��i��o�;��+e�6�&�}���䳑��)/$m�vM��4�6�3���F�m.T�"�(ww���ȇ��%�Z�K�7a�,�K d��
Y,�RD�Q�յ���?v㞕�0�	Cny�ʹXV4�I��K5�|�:�l��r_�ZGe
�"�<�B~���?���b���5�����S��?o��wb�A݈>Q� �D(��z!��5݋��v�>�����z!����;���.�E�(�{@ohl]���;�Z�*/Gi���ݶ������m���?�a�=ע�����{Xok�a��=ע>�Gވ��z#�D}菾V�����[g���m���?��z���l��D�2��}����?m����m{m���^�l��׶�?m����m{m���^�l����m���g����m�^??m�yx���������g����m�^??m�yx�����"�]���al!��E�l�v�=�]���al!��E�l�Q�ʰ�V�k�m|����g��߱�ߝ�l�]�U݄B��!�{�/�߻��%-'���J�U��0��r�nZOX�]�v�$�l����d2�[�nj�ɕ���o��ni
ێ�� ��u���U˞�;!W����8�������?�����/���'�܁�⸓���h��s����u�UFXAJ�eW�E&74����A3��+�=�)*�M��)~s����l�4vFH��\Yjt�Q�ʶ[���?�BA`�������Cs�s���-x�"E����U:�佖��?r���Fһ�{m��jP�P5�4�L�[��e���fh�%lK��nK�HTf䅑�v����FN����eu9�6�ǭ���-�w����^�:�:v�պ˛�bi�?�䇭�j5���~��O�����|+yy7��p洫u2k��e��ǆ��c?���&� �aR~(V$��+μ�3�VEm���
�&~��Z�!~Fr�)"�ە��,��0d�,�݈ܦ�}�u����:)R�b�+9e�~��6��ɹ��*��m+;�t�z8��z�{���c�^;��>:z��\��o���w����V�`��+|]���eo�����	[����K��-�`>-�z���h\@�T^9���?V�ag-T^9��e��x�Ik%@�㟩Y���o��R���J��q�z`��o�Kt9C��$:�QZ�d��E>=e�|��(�1���2_�%!vgr���,�K�n�Or��i�XY����/V��V�?0���z����AgrZ]��ʵZ�["��3~�%Al�^��ܽ6��ˏg%s��W��)�k6�:��D~_YmÝ�������u��T�*���J�n«z50�}������k;[JuƲ�an�J�N"���S7���&۬�ԤtWY���BJ.(��_��W;[�[�2�˟���A�v�;�]�Ʒ��G�)Kw��Jk>ʲJ
!\KqIJ����Yn,E�S��d�ǣ��Yg�{Z܌�vw��ׇm7>5�u$*Bߕ�4��ć!i[2�
�og�����$�m:���b!���|~O����q~jwl��(�^2��~!,�D��Z��D$L�%Z�t�'���2V��m�?���m�(B����6��@�c���z�T�P��(�C[�{�=l*z�T�����g�]�P'�]�P'�]��'�O�@�v ���{@l᭤5��������(��oh�5ʆ���������!G����i��2�~�*Wg���߽��{��>�Gދk�wc��}����ֶ>�����{z#�D^~�����>�E�菾Q��V��������G��[g�ߩ�]�jlkI;ѥe��wa��]݆��wv����k�wa��]݆��wv����k�wa��5膻�ע��^�k�z!��5膻�ע��^�k�z!�D5�O�z(�C^��ע�?D5�O�z(�C^���������[�4Չ嬸u��*!|!���������ܭv^�J�+6Xܗ�9�
F��e��Y���X���GY�V������ܵ'�HU���T��
��a�IR)J�cm߄�X�t��R��J��,��m&�$$e���v����E�=��#~U�&U�?r�^�qm��҄��Æ
�^�V��x1��Ս�N#n߳D,k�;�!�w|�p�䣻�̭�M@�⒢�t�?�2,h,��n��\��(�"�V7���pXсτ��v���vƁ(oy7��9R�����/����xn+}�V��N؄�B�B�T�����A��;[M��)��i�a�����)�<]ccն�An���g%Gi�rf˻����k+����)\R����H�K�)���(n:Ww�����!����69*ĕM��%&�J.�0���ůq��j�_V�\thڻw�m]K�O�,�Sa��ț�e�V��n�%�H;r�b3�^������[��E�Y���Y�ҭ�����2��<����Ӵ�a3~`���	�#H�+呟{0lp,?�vdI�l$U�V�}��㥨Ǹ�G֭�ȥ/��ó�UF���3���,�\�x�{�T�ZUO��9�ύ��ǾG␽����u/�b����[���d��Kp�>���Ed}2���$?u>����)"C�e-�je+yO�����Y����4v�\z11H�v��T�Y"C�d��lW{���c�^F�T��/O�S%�=�)��ҡ���VH�ì�,Gn�q���u���*��[�v�eR}X�p\���Y,��/WF{��9�e����'�X�+,��L������6A��)��]�}���w\D*��J�����~Wv�P�������%�?�vvP�M�]��bq]Z�jt��J�dr�]�1��W%���*��NP�B��(V��4�o���"�t���oyT��l��%l;kz���h��,�{h��K~'�vP�o*/$o-���=�l2�/n_�ݦ���'^�����r2U�p܅c��-����簅D�d���W�ԅc�{��2�\�M����ww?�b�2�Y��U��bMY��u�:�w�,]G%�ݹj�nV���;��M���R��dC;*�[��i>F�R�c��p�o��X�T����������@�BnoݠHP<��d*?/e�e��%-'v��P�J,�#����P����l6_{�~ǵ��|�k6��5;7�!wc��������g��B��S�
r�MdA��7�����elb�A�Z�G��*�:t��^!;>D6��Ǖ�5����[�c@|���~=wv>�����[kb�l]���4ƀ��8k[��.��g������c������o�������S
m,�2�^y)���罈7�� ��؃{@ob���7�� ��؃{@ob�ݠO�wh��]����v�>�5��7�� ��؃{@ob�A݈;�v ��؃�wb�A݈;�v ��؃�wb���>U�^�G�e��[g(B���o�)P%�X�B7[�ܿi��oڧj΁����r�q�m5�Oco{g
�.]�KV�!�=L��e)I������-x�~�6�R�H��U�ˉ@��b�*�-Y|�;��b�����ϳ�D��U�����N_�j�M/O�[u�$�������������w�~����і���:�'�O�8��$-(�v
Y.���W�Zȍ�lqv6]�-M���\�2������%Y�U�i[��������J����L��+�����6u��+M��V�q�Qےg&�W'��^O#I�}O[��d����Z=��Ҥ���KWX��վ!c	���o��7�a��4\if�d��u�!�݆�i)��x����w}��b/��:=�9hU�+�;�e��+:�+/��r����-_Ů�h��6
�YIN���洣zk�ݫ��Wo�����	g�����gI�����e]��+�6�*��"6�7Z�BB���v[;Y��^�wMr�6��ܖ�Z��ۯ,���S=�D�/a	��2Uc	*�����Bh�!V��}�O��br�X�%��4V)��nr:)������m�9Y���V�J�I��������$tv�\H�ݮN����Ze+y���;����Ҫx�v�\Gk��j[�=��vR�ƦR�������D����*�>�Z��}���������`���Ǫ\t�C�h0��=R�iu�s�t��?C�J�}N����+T^R� ܏�$|��m~#��n+��;ʬk�`����Y\���MyV��jѾ��v���G��dO\�7��>/+�����#�9Y*�S!W�e)f'��A���T7~/wcJ��C��݆��ʲ��gd�U����/����u�}d������|�&Ki����m���y[�6�Sm���ڒ�tH?��݆v˱�iV��Y����jd���C}��~W{�X����m�$*Ɲ���viJ\;{:v���*��0$�V�?iA�gq:��m�_v�%X�G�)#�F��΢!r��gpc5�%b&�BOa��+=s�5t�m٤H�o$�c�r��c�(n#�[���*�M��ǳ�i/��ǳ��E�S�@��}jT��~��c�;܍+�P��H0�Kl'nR�������å��~
�%`��k��-�+@��~v2rTf·�c���2���<_�moG*/k
���enM�v/�U�o�;�N�
���f�������g��~6������e��D'��O{
kaM�A��61����h�66	C���17<��۫N�`S��\�?�cm���5���~z��z"��]݋��v�.����l�1� ��Jg@la���g���cm(l6{l����a���������?>U�{T�1�=�A��OclaS��T�1�=�A��OclaS��8��:g�g@l����B����OclaS��T�1�=�*z�T����aS�§��O[
��=l*z�T����aS�§��O[
��=l)�����ƀ�D��w�y�UG伅�=���#���F����@��i5�����z�P>��=�nXh�b~����YK�+�M�%Q��~����	f�L��X�qE�++�����3F�#"Q��;;Z��b�T��,�FK�as����&��`����ӵt��hJ���0���.<��Q�"��������xݻv�M�k#՝�{/����°9�B\o��I���Q�{�%]�̊�O�U���Yy5d�moe���AAF��쓴���<�!���V䷒�)�}���Cc!F�d+�K./"?[��[�;�7��B���u��򖬋�'�o���t�Z5����Kr/���3K��7K%���)��D�@���e�jݪ��dB^C����2}�o��?��%��B� ��T�6�%������K�~�\כ*�.��u2��ڻw�����Bh�a����4g�6�����r/@܏�坻�u�:h�?�@��Y,�K���ev��]��+[����.5y6��m�[{,�������~+;�,dd�[�����C��x�VVe)UčO�C��,������z^�Q�ǯ���������;��KӨ�s��x5��q��NIk'=pbKY<^���4�-�}�?�-t��B� 8[������x�1녜|�$���r������^���v�Ė�\�^5q��H��y��󎗧�A�_�GA��5@��%d1++��8�������m�vRC�e�=��v±ݬoܿ0h�V����(�
��.-~V�;�'�Q/�9Ѿto����z��x�U�y>mͺMn^A��k�V�ӕ�#j"��V�+S*�by!���/g��d��V/�6/�S%X�1q�����7�v^�[o;l+C~��Xۿ+rl�g��d�Ju]m7Fǆԡ٣e��H���[;L�+��Xlc��쥫e�I�.2��~M\w,z�%�;�O�'��ݰ���������"�P6����5�m)~_(~Q��W٠�bcr���d�%Aj{-E���!)�6�7�|���T��Yʫ�
�����|��|�.�/"���dڈ��im�+1���gwr�Y���Ȃ��Ȍ�Ro�,��}�����zu:
咖`�b;>,m��:�~A��z;d/������'����Cml�evNJ���`�2�N^P��������(��JVB�jw糠a��0���k8�M�϶{>���g��l�g��m;g���w�y�Si���6����B�HSg���3ջ,Z�Ý��9k�";��2��n��)p�塶�Q{[*�^������������[:g@l��Ȅ�P��"�D/�P/�D/�P/�~50�+�Oi��@�i�g@{aOlA�7�Ӷ{O�Ӷ{O�Ӷ{O�Ӷ{O�Ӷ{O�Ӷ{O�Ӷ{O�Ӷ{O��=�*{T�0��aS�§��Oc
����m?O����m?O����l�g��l�g��l�g��l�g��l�g��l�g��l�g��km��Y]Ʀ���%�����X���pY.��v�}��{�T�R��x����e��Z�˔^����7�4�*�v��d��6w�!o�5lw,3rH���V�B�H8��/	_r�'�Z׈D��d�m�<�5�ɿ,#�������I�yʫ��h�䳸ܤRK艫�1u�̺]j�^M��U��Y��
�8��1���we)V�R��g&��g�w��U�cf�H���dU��͌�q�&�
�a��/�qq�����K+ﹰ�Z�ݖJ��e-�YWe��i)��{ͽ�f�e���:l��(b7!��:m�JM�A�I�҇���ݬY�G��VYT�g@��3��,r��|~�v"��Z��a�Ձ��E�+:����*���p��?�}�l��M�ʈh�� u2��c���	CY[�嬹_��aS��ݦ�VP��~3ah�a*������W���y��G7\|���a�E�g���@����������nV�
�����!�Ȃ�V5qyj�m���;!��N�-(Fɫ���̏�����8L�(n�����#"�O�Cw�������Pm>+�|���uO9��Z�����s�x5/wG��r?��~)�}ss�x1�Y���J�K���8C������Ix6�}?�?�y��o8���,�|BȥK���$u*���cؤ{�E*],�A�ru�>���q������8UO�S>$h��������;���Z̥f;�-�+���R�ۮrE����"��������i��+��_��ą�e��{a��-�_��4�%K#,h�F�٨ޫD�z�﯍�ϳ���z��2�Wќ�1I���la]ܽ��)`V,�9|�7Y��ۦڠd��{=�b��n���릏��[�q|W�*��e�4�OD�,��|�w(T����-N���Z����ns�ӻ-��T��!������U��/K����������%V��������_G&Wc)g}�_gX�JZ��މKv�Wn<�S
��������[�H9L�b+�խJR)��M*�����%�:ە~�rԕ&��a[�I*�Q��-"�(Iݾ[~e�H�~[�B�Zl]Og#x��w�o�0m�VVO����M,�E1p�|_?[���ׅKu��g&��We��:'-�_��ғd�����l�ir����i,1=��<��[�-�?D_������/�gN睦��+}d*�9B?�Rᣒ�d�M7m�J�B_S��j�\7�[.˅��l�[.����i�Z��˵��k?��˵��h���Y*ܻjʩ��,�R)[�]��6�?r����{d�ݝ7��welb���61� �§���e
�S�=L)�����B��D'ʈ]�P/�v�ߌ�k-���OY�*!wg�aj(��5�7�;Z����g��ֳ��gkY�~����Y��p߬�k8o�v�_��~O��>W��_��~O��>W����gkY��v���gkY��v�\-�e�~˅��e��p߲�l�o�p�\7�[.�\-��.[}��l�W{�}؇=f�T�I�e�b��E^�Rqe�x�kn#ǷCqZ���r=��Kyj�qJ�Hꝝ�h�I�u1�6|R�$�
ܔ!���/�lC��[����X�-nF����2+u�zO:���__+���I���6R*o"'�n���G�{#������4��Zy�7V&��Irۂ���'�Z롇2��-l�_%C]L�S3�&<18���<EoA�D�`�����*�rc�J�r{I=6�_"�G�'_a(j�4�yQ{n.'M�=��^��wn����׫��׳o�B�"�V�s��o������V����O�@�F�d�|�*���C�Ym��V���ߤ��pyZȾ�-���!k��6��aTrq
>���]��؇=�n�T^M��$�}6�/��l��,�7S%iD8k4���m�d>���*w	��3%漼��U�r��`tBh���>M�ő"ݳ�p�Y�����RU2��������0؃�g�Y[��h�C�c!B���&���E*R/+c_	���>��>6��

3�&���ҡ�ج1Y��^V^����,���ej[�$��#Gv��"���A�h�ֳO��k0�n��Tr�K��' �l�Җv������{f��A��a��G[���11Mn���64?g��Y�f[c!��p
e+yL�o+4�\�!���9Y���)��qn��5?���q���-��]D��Vm�������?���$t�� ǫ�+%n^���$���⒬�X1��(ɷi0xeMw�{dŖ3�M��£uFk��}���@��"�}���٫��J|���b�,dۼ�!_u�xm*+��E��hxv�)��a���J�!�!�qu�͜�a���obd,�~�ʋ��d)?���+��B��B��
2�:�.��r_��Ao��55��$�X�H<8;��+r&P��݌�V�e�U���Y�m#�ج���$=��F��l��)o[�����&iKWn_'(W�?9��nܵsV$�-5+�@�b,}�O�lm2a$Cy�u�+1�"/�)@���ۗK$W�dڜ��Y�Ղ��D��u�mk+���)ؚ�ݻ�Ǣ!X��i$)>����϶��h�*m~�&���Ӯ\�-��"��.Yx�iKOM�rJR��Id~&'e���V3@��D"�%�����m�)\�.F[��w�
���݆���e62�l�(oݧk�vW�|�T�ҁkS�~�~z���w��ߞ�~z���w��M��v�]���-��~5��KI��)Ctr~c����2���+N��4\�/������Q�,쟕M���Y.F��B��S���~O��>Wm�Omܷ�n֛�����s���B��W�.�X��8X��YhU�B�!w�@��!w�@��ߞ�~z���w�ߞ�~z���w�ߞ�~z���w�ߞ�~z���w�ߞ����jxZ�����jxZ�����jxZ�����jx\�����ߟ+~|�����ߟ+~|�����ߟ+~|�����ߟ+~yk�i
���c��խʐ�RA��YӢ{���d����,�HZQ:m�-E��ǅ��(k��$
��X�9)Z�J�t���w%���X�hnZS߹Bd�����GZ�K�/����w���w�z<>�\�A���� ^h��2϶,�*�|+����d�����M�q8�K9�n��`���_r�륑����g���J��հ����ܥ���[���h�n�ՖZ����՝7?�^��[
��c���r2T�d��퉱�ө+2ݍbM���|��U�������u��K>!��)iv�����;���j���W/Fҷ��p�a���^U@���v�!9) ����oZ�&�$M|��|�D�(m�)CM�a������Q�RR����i�W)(I��x/FK#c����!R��?#Ek<�F�%��i����2��)�Q{n�/���Q(ڸ�w�(��XtU�j����O0�Ϲ��=��;y��G��-��m6?�[q���l�[��b�yVYKђ��7$+vU	��B��RDv��퍌M�~���|��g��_&���G��o��Ea��NVe�϶�\e"�:�A�"�x1#�x�=��/�}s��mq#��_��g<Ϗ��p��,A��>VqޯԬ�B�>Z���'�����z86I�z��ϽP��-�{�|��w�����Y��:^�G�0osO���/O���]"� �pĖ��ĵ��2O�\п~���C0��������
��+��9ꖢ�F-Ӯ�,���q�������g�k�$��ҵ�ݔ"����x�X����q�Q��z�yu����r�<&��'W�˲6J��E麲mϹ�O�^����l�?.Tt�r�m�k%����������I
�u䓥-z�;-~�/�J�ô�}�p��lG�TRU���R�@�2W&ҷa
���5����+��>t��67M���ܾ$�b;[�)���[�j$(nv�,�i;l�?n�;��Ⱦ吔�Y�
n�Z����N䡹٬�D�[�u���쵌zB����m�܋fK>)����^j\�(cgV����v��_sB��q
M)˟Y�ܲ���3��14�JR�¾��Xd�%��x��պI4B'����?����w�V�C�۫��攰>��6�Y����?l�ZU���(FZ�p����9�]�U!\���W�rW$���w�wQ��gc���Y��Q�T7cqX�ew��E�ey'�䞛���e�nF[���b8g�ឧ���b;Y^�W���{i�(n;m�x�=�n��H�Y�$�|���96�C3Yc�i�����K���g{Y��w��ߞw~y�����8g��#�zn��ݷ�.�.�.�u1
�n�����<���g��c��p���7$�ܓ�rOM�=7$�ܓ�rOM�=7$�ܓ�rOM�=7$�ܓ�rOM����S�=N��;����S�=N��;��r2܌�#-��r2܌�#-��r5��g#Y��r5��g#Y��r5��g#Y��r5��g#e��\��ۻ��Q�v]�׻�����mJ���	�q��Ԫ�XҁRO5��7%}�/nO�ŵ��i/�٭�j2��~N˿�ȵ���M+?����VR�m�Rh�������86t���DJ!*���#1|(B�5'�MɃ_�g�ۂ��iF09�u�ܯ��Wщ�F��N}ōzO��ǃgk6��b�p���e��זZ���竷"����6�d�����'��U	�X�uہ���>62�&�o��x�3�)�,�7�:��JM���%/�喏孱��+"�_X��ܱx8��6BܧSwkr���7!��ն���ݲ�#�%)o�56���˲��\�Nwa��i�i+�m��a�����O����[�<��#��~_{XǱ����+���y�D ��9JP�1��ݽ�g[M�IY-����\Kud~�!vqp���ўj)~v�ї���ڻW�/_.�q��
�.��5�D��!Ce���(E�1;�~vS��}�mc?-���j5��^ݜ���e���}&EoM��鵑�)U����~nqv��P;7!��4ͅk�㤵.G�5����H�������ed�S���w/��?<�����r��1%��sB���&V�����E����osO�z9G��;�sB�z��s�eo����4*��}?>����}/G(�/Oy���R��Ƒ�����~��T�P:�K��*Ck��ipĖ��w���㒳��W;ٵ���F�P�|�8د/��d������b�ͺ���R�u�<��ӫp1�2��J��+����X��h���:ˏ���X��wn΍���/Z�|���y���rc_���[yl���Y�b�e:�c���[.J>�njo]��o�T��c��(W�1rz�C̅��Q%Y�9Z�������V�c��7�uM��`b>Y+l����N���i��>V��c���������R��d��:�^)R��1��#���k�i�{:t���$��j�9�ǳ��.J�G�W�]��r���ݏ�/M��l���?S�����;7��Yv;�	Z�g����a�a����頠�O��-�,��7�؇�Z�"E!�`���8n)�V�'M���~AFl���.T�n�<�*����&�����o�'��������e"��V�~&��k+1�c�'����T�J�W�.?8��!�w��J�\��P�JW$��9Kn����#n^P�f�+}t�&"���a��N�rJs��'��W�znI�'�䞛���i�nF[}��exR�jR�I\+.�ۀ���䤩6/a���H\98��6O	�Gn����a�۫
ۜ~䒢�{X��#���gw�߿�w�~W}��#�x��o�vߦ�;�wgXѲ���B��8g%r2��7m��˺�����gxV]��{�/��OM�~[nym��'�䞛�znI�y'�䜕�9K~rW$�܌�#-��r4܍7#M��r2܌�#-��r2܍7#M��r2܌�#Y�<�#Y�<�#Y�<�#Y�<�#Y�<�#Y�<�#Y�=���<Mf��/��Fe�ڲ��^���gm�u��,�U�ÎE��%v�¤X���ܤ�;�w�V{	J�Q%iV���d��T�K1鸬=��&��oK;(K2�^�Ow�nU)D,"��t�����?$�$�G�/$��(@�7R~|�!"r#/�¸�v��P�{dn[����h-#29ʳ�`H���j
5}U�k�\�1����*ݖj���~J��ፓ@�iX\pʒ/�d�d�+:����r�1ʬ�0�z��״�V&�VE�a�³k;Yr$.�K�!��ҬW��ǃ��߂�ׁ�Y�ȁܔ78�0�]7����Ww����f�|o䛇��)~o��7�|��o����rۙ�_�5��r������U�]�������Z/�˷��s�^�JR���e(��m��2x�N�/L��m������v/�N;��Q���r�Wq��qj����Ӫ](���qdju��gg�%[r���'ks��񴎾R�6�/n�sі�r�,th��^�&���6��o�d���Ë_VYI���*��\��(5:���x�U�G�+U*|��[�]��\[�Pc�Z�J��)s�Ed|:��mk�-���0;]�)���2���S>>Y8�' ��#ތLR�-�˟�O���u�<���)[�L�R���yKwa#C����#��e��N�[��#ތLS{��kv=FR����{�x�R�H�ݮ&�K��j[=E{�����>簭C�{�ʙ�ۮ{-��/���$��>�]���%�)c,��:���}�����qQ�D�v��z7᪽�E^��Z�W��rJ�}�,�-f�/�u�-�knwr?%iCi���眖���xC��*�!������b���|���dm'&��l���F�o�U�J���V�!���ì��l����Gcn/�HQ���Y�JT��#����v_v9.�� ��5?Z삔>2r�Sa��؊ַW-X��r��Eg�J�e��w-HQ�,�~��e��]���l��*J��d�(�k�r�$�I*YR�)ٛ�`�$a�|L�e��mӒ(
��Ĳ�+H�%�Y��Vb��%6F��#�5w0�+����k�wkr>F�e)���n���P(�m6�%s�d$�4n^!�J�@��u��9�I�ݎ儡,���[tҭ��͝�X�H?�i���\�C�(n�Z�o�w/��.Z�yS�I
ۻN�f��%�R��D�Ȕ9-�KnrU�rU�zm���s�r2܌_
����-����/�}n������\7-N��&���@��z!Ym�B?)I���;|4v���²�|,^��-��\��\��\��y'��b8g��#�zn��ݷ�;o�V��k�9.�[i+m�߿-�~ˆ��-�~��
����V6���se�Tu����]7J�J[�+m�߿+�G�v?ȏ�5��r�ICI!j�ĕ�<F��V�;���;mN�;Ȓ�-�K���b6�۔�l��x��v�<F�-�~��ym��ܓ�mߦ�[n������r�L^�R�u��r*܃����J��#j㉻W���s�B��ȼ���'��8�LΦ����Vd��T�y��%*�D�K���ܶy�}�I4�Y_�*䒢��;.�'M����P)gU�o��%�З���/ap�Q`�AP!Q0�z1~+X2t"��#���_r#G����-0������-Q��M�>�e%�5\9�������2 wl4g��dD�e����og��@�l�r��W�i�����Sg)D�f�J�\�<�x�w<�%�>6U�"�M�F�:�~B���њ1r�
��t�ܖZ��P�R��z$����#���/������@�BJ�<�e���y�kڧ�v���W'�m:Y��ijqy��٩�P>\�.�g���)���e�ov9mn��J��5ϲ�z�i;'��Q]�s����וn�ќ���gF��L�}��3��k�8�n�����r��9B?�!�'���M	᯲Ӛ�\�K+!�;�Z|��=V��-���q4��./_��WOq��o�J���ʃ�*j߼�[�}>���a�=��*?,v�+2���H��U9��d|�o�E`R��Ht9YO����/��ǱK|{��3��S8�Ps��+"����B��[���/���x�R�C��~�G������mc�Y/�p4|,�T�����?깊�8�?k�í���%�ڟǏ���4����{�P*p��H���ik��|z2��N�[�ǡ���l�w����D1NKԫR�i�%6B��wE:0���WSN^�����g�(��R(��V!�aۓ�1���4���7Y���7��'8������5��R�����A��+�1Q���{�U|��ԡ������%ou)P9��չB�wc�k~��*F���ʢs�}���ݒ����E��E-�e���J���D�u5�y*�R�R��� ���T�H�GQ���eN.U���J��S�(m��⫟m�ݐ�+:W/!id��nQ�/�ȷ�W���F�����NA���jV_������݄W�B�a16�,�B��Uŵ�I��U3o~Gu0Kk���i���lMKec�ܨ:���vU]��Kx�4�l��M\�!+r}݄_�:��/"��8���J���r�
՜��/M�b"�4���7i��+I�ܻۻŸ��J�K�XH�m{��b/	e���³H=�aZ�B�R�a�v��"�RJܗ��Q�`��y�/�����v*E�qӲ�*�N!_e�yK�)!�|�Z��ǹ ��M;��6:Vtu��=�
�r�v�2T�9k,o~�_]%o��R�(�]X�i�n�y' �}�c�7�{g�����U�w[*lE�y���]��b;�t�����\�)p��]V��G+�~�����|����X�ărV9�D�����B�Js�B��b��X��v��ܚ��#m%r%D�Ȓ�؋��)�.S�\���Or�"�<E�x���)�.S�\���Or�#m��b6�W%��:�*~��YG�����
2�%�ь1��VM���0/�Q���#�}����Vmf�ZěB�ۑh�F9�XİlO������;^j�K Q�Q��o8w%�eƌ�+
F�&��h��W�ݸ�ooZv�黕wl�`c���	a�6��$��Lm�p)�O��bh���hɿ%�r9�m�Y�pR�64	do��gVϚ�Խ�U�<��-x��ɯ��a��:�R�.A�l�^e
��Mov������n��d(�������H2}\�&�?^�G������!�mܫv[C��gm�1~��/�_r�^]�*�)Sp2��A�y�ra�y3d�n9]�t�W�|�V����Ht�D�O�z>Y[lC���ɒ��aQ��TB�H�j�ߑ�K���0$Y���;�����V�;��,4Un�ݻF�����^���_�0��������\\�C�v��ebX��$���.�F��J�ܴ���Dn�����m:�_'�����ߐk�-^-]zJI5���Q$E$�ܑг�+<~��K��=�l���;Ǌ|T?깮1N�,�㐳��T	-d�}Qg�ި^sB��/O��h\���t�or���?���W�����#����7�|ܯ�������ZS��u�܋2?8���(�V�$/�j��pVx�:��q�_O�a��o�p�wl����*r>�K�J���"���\tu,VVԱY[�T�K�{c�ݧ��v���۲pȭ�#`l��K,���~d��ᴼ�^�\6��tf�F}Ȥ�ݓ�E��1}�V���E�V?�qv��H9��<O�t�ge����v}�m��k93�1Ջ�g�i(��n�U[����n�K�o�t+��n��&BÊ���ߔ�[���I/e�����7ʍn�'��񵯓S@ȏj7d<�������4�R����yiӬ�r�]7�R��t:Sm�j2]����O=��^{y�V�ŗ�Y�b-��nPݝ6���[�T�����^���+���1�q�
��d�]sds��vnl����.UZ��e��kw~č�_�{hZ�aZ�]��7�X�y\�|����
F��	2R�}��[��l�#����&�m�������q�J���a��.Y����{z(��r��BP��%*t;r��o��/��F/����s۹a�j���N��4�j��`rU�����q��|�l�?���ܱ��W��9�޹[�\�7�6�sq)p���������r�B�qa�������9���&�_�����IV|9܍�ln����*���a�����U�7+M����k!�}�)K]���%~K����&K��V��ض�sJRU&��|�ێˤ�G�5�x}�=*lG�w/r��z��)�Wr\Tq{�-��n�7n�6�~/u��ewRV�J�NR�˺��Q��-J_��|2����ح�\L�M��ܙ[�%rb�ҕɒ�ex�^&W���ex�^&W���ex�^&W���ex�^&W���d��V����/@ݿs�,J���%|OWW>��Y��#���mȞ���h+K��_Q��/�m�5��x)�aAsW�2%�4"��ɳ��B��ln |˼�u9�o��,sa�v�~aՌ���M��_�JY��"�Ce��������X8a%�u�����������c.���~�ON�ͫ��E�f�g].��7�/����τ����Փoȿ�F����Bf�.����,�~�j��k{��E�ʝ۔�3�Z��AB�c)��2��A�ה0h��mf��#b��e_�2j��k$g�hn<��g;;��/��e������p�%.y�W�Cs*�	�Ḑ�*�u��a��ܮ�+�)S�)�M��~���m6�Y��i��w����>P=|��=4UÅyV���ڪ���z��:5n��V�~�>p��QQ���([z��4O^�6��,ѿ`����
�=̍�+�dQ0���yUĚ�{��)|�.ѵ&���p$�v;��V62(T7%��Y��G�����~��g�����#�H_9�8�K��|��x1��elG��d�Y<<i/�><%��W=p���H�x6��)���)���+<~��G{�^��IiO�����@��<w���+n{�_��+jPĖ���7���iu����+a��^����+�>�]���-�3��G�☥j�\Tj\uθ����>�K���v)Z���n�$E!��1+5����@��;d�μ�VA��6;.K,����E���^U/_��ֿ������ɫ��#8�Ԓ��*UN���eYܯm�J��ܭɷ�H�:B��2�_�܈V�V�%dJ��P+����/�4�u$�m����:N�.��� �)5s��D���V�F�rd�laV�j�%[�����}��e�gM���Y+m�e��~�Z �w�X���J;�ݷ�l>R��v��Q��$>T_����Yl$m�*;��Ya�}���Y+�Y$i�$�mƣ�?��4X\�-WނZ�vW���̜�R!gn���Z_� lx��h��$_K�7I��TR=N|nˊ�	g9F�����v����R&���h�L6��v[�)f���bO�����+|�Ԝ�ԙ�	?Z����9����y4��ܳb�+<�2���ʻ3�qh�ܴ~[bv\�;ѷ��/�v��?��4bO'm���Ѳ���K%c���qv]�ϻ��d_�,��p���6�A���I[���+X�Z��gd�'�
�����h�'w^U��g� ��1���չf���ٟ}v�v�׻ݣ�عg��W�?4|�V���wv^J�ш��V�4~j��Td�p�ʼ<�m��J����ŎA�NRϣ��c��Z��3Ya���mN�l�$�N�+��˷V/��n94�՗n���[�_;r���9��f�v$��;/m�w��uoU(n�)nNRܜ��9Krr�Pܜ�Ĕ�V�J�I[�+q%n$�ĕ���V�J�I[�+q%n$�ĥ���1{�Kn�/���u�G�o�na����_�'\�Z.]��2:���������櫭Յ�EqN����>�u�6��/�^Ee�W�m�:u���i�,xdPQ���1�c�P����Y�,NL��Y���Ȃ�*�NՓb�k�Vw(V}˒KJ���,���X�f��w5�l�w}X�Y�j�yI�nwi��*�]n��F�Q:_�Xџ��>�2+���\R�E�_���˻q�&�V��V^�-wmզ�+{<�Z��ȧo��(T����V���ܔ���jy#"��.L7f��2zĞJ��Zj�o�XX/����@#2\�e�{�w!%��8n��;����v]�v]�}L+϶�a�۵N�S����]�"�.�	��v�����[��5��s���g�R���3�X?��v�ڵh㴙/V��5Z3�UV��iޫ/GkV�4N��[Xla4��	�ݰ�b�θu��	e�M���rk�D�hb*:R(N���эv�e%�=60Q���5~�~��e��[����aҖZݒ��q�v��J�ok�?m�ݨ鶒ާ{]���M��r��^v�N����)jkZm�����)Җ�ۋ�E�(�o{�}�KQ��I��G;���6R�{S�d�?e�m>T:nJ�m���y�N�16\�RA��jܥ��J�-Z�l�U���X�d䭍+-�䶖���e�H��췲��rދ~Wgn��e��&���E+{L����8e,�f�G94l}�f�D_i���9}zul�à�ڵTK˫���Ǉ�Ɖe}�D�M"���RAV73���)~U���H��Cѭ��)ҭ6ǶA�ȸb��xd�@��;b����N��b�:[,B7%���]��93���2���k%����ˏ�JnWJ�ʹ}���aٖ����=���B�ɫ9k��XYg�7��o�#j{5�߲V��E�4��c����v�i~S3��SM�%(��n�~��"ԃ��*�&��[��52��U-�S�\�>5��},5uq��n���2Em��[�~s`��Z��D��Fhύ�,`cB���R.u����j�2����
�Jϖƥ@�ܫ�ό��Ar�xĪ����96���C�Ags�U�j��B�n[k��>�c�̶�i���5��W�R�v���|Ȓl��-[V������K�e[>--�ܕ!������m�T�~�����[���5:�-�}�u:m�mb�Kv_���%��K���V셯/�"dYd�/o�M�,�nɪr�N˫��ہ�ȫ��j��߁�7lU��lC�$C���%ʌ��W-�wM*l�r�26R���b�wp[���d��~'r�������1~�]�JU�`�h_��O�,�R���$)6!�j���S����Uw��.��$��ԅ���Y�{ud�oU�Sb�5���l7��C�q�IM�!nє7o�7o�7o�7o�7'(n�)nNRܜ��9Krr���-��[���')nNP�J�Cu(n�ԡ��7R��A�H=��e�H\IJ��\��We-��r��v5����V���]be�D��I�ԋ��8Hl�__��)�<�q�	�v04ul`��?)
�n�`r�W��Mx���0 kP�W$}���ca�##�
�Q�V_�X��:�U��R��)<����ww��%-�a�^�l�e�H˰�9����U׷a(igaWɳZ�h}0��Z�'�W��p`n%^|�RWӵh��).�ް�_���D3��n�%���rY$��^?�g������ѻ��o�h�gn[�>˥���2?��Sq2&�!���dcgnR*�����#Jv�6��!�ʹH:�̶w_+X��kՔ7mwk��L2����0��Yuj�xc2�TB����+t�eg)#���!�r��A���͆�O�K��ToL��%%��T͚r�gF���ݝYz6�c��j�\�k�?r�edRU6_�Ua�,�X�U���@�J�������<�\K�4nJV]��_�df~�$�O�K:�+��Og���$�T?;����_l������ֳZ���Py"C�Wm�:+�e�)#K�[�z2�<Lє�����DS/O��+�?є��|�:ϕe��luN�s������q]�g����Kp�>+#�����/l���{eK��ǱKuFK�t9YJ��9Iݓ��r��� �k��;Q�m2��E�ko�pͯ�s�%mθ������� ��9k��R��u2�\S.uƦ���;n�;�
�s�FXv��HQ���i�@����̞֨˗Iv�WmK��V


M'��,i$Q��})�rJ���=��C����D"�D��ʦ�Yy-v�]�2ҫ��nl�2�N��pܼ��я�c��BJ,6\V]��,�~+X��E�#g[����r���w��TWe�HW.T�M�wi+�ỷ*~�̥�GV�O݈l�q}FW_�����[l�¬8�2T�e��S��m\�&�7J����≏�%�xT�R�P5?G*�ʯ�q\S!���+l���������'o�)r�#�����̷[Cz�K	�ό�nY���\'a/'�J�~F���-�ݕ+�շ�l���5����
�D3$�2���6���n��Ȯ2X.,n�4�q��X�ȶ�!U�Uo�� �k��^��J��v<61��9Ws#;�*�nRb�T!!3���>[r?��r#�pRz�*��h&�~k-bO��rD!-�����E�-6�S�����'e�)g+e���:nC%rǿ���/S�oǴ��Rl������ȈA\�.$�h�F������W%*�'�J�X�t�}�T�EN����V�q��z���~2�N���+=�,p���e6;n���f�۪y�=+����B��!��m](Vh�6&�m���"7%����I��G���B��l������I~-'C�r�n<�ZU!b�(�{y땚����kk�^˶^˶^˶^˶^˸�����;'(vNP�J�Cu(n�ԡ��7X��/���b���/���HZ�J军�v����1}���R�YeL^BJ�Bң�`פ���4��>d�.K�3��\�V7گ���g�"��E����r
��Gr>?��Nݯ���[����J��bk���X�m4�l.$]���14��%�����8zʵsRRK����x�㍰�a����_��n5����쉌ⱄ��_��e[^W��g�Ə�nnKmr�v}����³听�Mx�I>��"��ɨ�9�эܓK!��TW�~/_�M��Mդ��q"����,��ɷ$-x���e�bj.δv_���ʕ���ݏ����:ݹg睸�$����f���!vU����!�3��;U���!�Y
��nW�k�\����2����27w?#wK?��x�-/-Us��V��3!}�7Wf��}�ݗ�G��ᄁZ���_O��U��ܽ�)6"BY���J�����?0�٬"zܴ���RO���� �5�Ri7XO�n?��RABBk��y�I��I:|:�(|�y�#�]�����gP:@�p>z�r��;��d�Ƕ��~+��J�>+�8�}���a�tS�����N�-��Q�d��+o�p0�w/ ����?���:�R�a���b��+�����b�ύ%�ݮ+��J����ʗK��
\��b���R���s��{��<����jP�)��rr�A���d�����mj���@7�4S�Y��{�4�˒����*�ېk��q7)Tg�}��&�B��cƫGG<�h�˧U��:�%�o��ƾ�M'��I咫���>M&�ǟ��`o���!��,�R�ѹ��S��)�z��{u�}���mnM۷�VMv��R݄���k$,�lB3��ȫ!k��o�E�~�+t��Z��t�d�B�K$.�3[[�|�d��䍬��P(�����'�6��\���LL���#JP������_6���)J!ɷg���"��~.�$���b���iv�
��W{��AF��3��4�ܽ2۹+12z��6R��A)Ƞp4�������(k�b7 s�j��&B��(|덛a������H0Q��T��ێ�c��%��;g��B�զ�Rlw')K):A�͝҉�F��i0l����O�4&�|����n��M��]��Tw�t=oe+M�-�vR�����5�h�ˇMÃ���r��*�M�H���Gg'��߼4,��/<�M�e������64��N�ҞJ?�M���o��k5�z���_���;*���Y�kK_4��6OL�|���kM��J�d�������"ߣ��ҕ2R��:R�qC�kv�Y���T��ɿ�U��?)J�d)�;��O�11|�7�H�k�r(��g�ٹ���Sm���+7o�����@�}۠u��,�Y��ݬy�ed��<\���۸�}�o�>�,���ϐun��n��n���uo��ߋ�HZ�]!k�-t������B�YuV]U�Ue�YuV]U�Ue�Y{.�ug �$T���k�$�����۔��r�X�ǹ_G"Ƭ�O�M"�ݭ��҂�҉�'�F6��f�:�-f�ό����v�U���s�b@��Lq��Q�Q�e�m<�i��1�tm����ar�I��Q���y��a03�nv����'F�վ��&=p��/�6�X�݄a�<Ԓ������v:Q�U��d��� ��`�ς�۰���b���Ky$\�{ML���j3�Q}y|���ݱ�{ca-�s�.����w�k)5cso�X��t����*���\1����,ᰄҁ����w�7,���D)6P�VN�*����F�B�Y��P5�RW��A��97tD3�e�PZm�ym��Y.R죩��IQ8W��N�Yqr�؛�.�1?���jU��/q�u�Oa_��F�5��ӝ�g}�ݣ}�n�V����Z��q�M_a���gaY}�f�S"�JP��~������/c�r��Nr����^V�O����߱�x�5�zJ���?g��uZܕ����������3�bVB�/G(�>zVqީY�z��S�s�Io�⹮8W���g�݊{��-o�p2{8��mJG����K����⹀o:;��Kq�g����YJ��0��Ix6Gt�8Y��81�3�~��ԿR����:��Va�)O�����T`��������121���6r4:�C�m�LR;�ډy���%-�v�)|�c��V/-����鵛r�����9���˲h�.M��}������}�V�^���?:'j���i%�{9F�3��Tn��F���[t	6˟��djeog�����g�qɰ߆�r�N��Պ��l���6}���e�̊M|*�&�l�k����w�ӅI��,�[nQ��w�~Jݰ�I�Z��6����l1Q�C�6E���Q�OO{����;�����_�ׯ��΁�ïq�[��WwvM!D9!Z�7-����(v�����򭽔+)N���;!ژ/�j��:ήKU�GY�'��Q49B!P-���֗��)r]׆Y�/���ͩ�`�Cld\Wn�}����J��[��(��G<�9���lnN)v#J[�ʭ����/�NB��+�<\~�2_"���H;��C����`���Xֲ�RˬwMO��e$(l_;%D(;;m+S�ʈK8l?����Y��ℶ�9���x�a��;��]�OfD�&���܋�r[a;8q�k4lg'+W~�X��[`��̼*2��"�"^�ƽF�WJ�B�K)ѵ���_�{hl�*��@¥�6�1�������]���do�R|
�&�S٩�075h����Iњ�ѱa�B�69Y<6�X�le�Vۈ�:�b�e�JY)V�����~&� ���)feI|�r��v�jw�ܴ�������P!�a[x�����2����;m�Aջ[ջX׻X׻[׾A׾BվBվB�HZ�]!k�-t������A�H:II �$$���t�z/&S�R��d�]��c�w;�WMɆ��|"�W5�Ej�%"����	�@��~G%~���
�
|�Ќ����ۅ�WX��9��y�s�����Rs�������&��vD��������_�c�s����܄����M�K5���K3���h���%!��s.�~+	?e�_,=P1�a,sFY���u�������i�����l�b��M��,��֬jY���_���K?r�BϮ�~�V?�"��J��SN�[t�Z��~ܳ��4�o�ո섄��_E���_�S��B�2[��k���z��*dCw�r��ip�r#�E:�&��2WN�!�+�vJ�k6��[z?23rk��἟��ڸp�R��������O'����+Ud��QFJ��y|��w�Ѿ�[�պ�uFj3��<��<ѿcc���&�]��[�s��u�Ǉ̚Og&�	,�����"s�r��嚺�k��"lq���
��_�ű�ҵ۞�ݵ����+�C��#�I�L�o9[�졦�gvr�����|�?k���z~�i��m2����+!e�V\�%m$:n#)M�e4�������a�n�NR�[�y{f[[o�Va�
gƛc!�w���&)���{�LSe��UN��m��5y$����%���hy�EFB�Gd-dw���[;~W{o��.|�E�cY�lk0V�٩����+}��Lߔ��>�$6��%g|��հ�c��N�D��c��ה$�k��e��6�WZ#:�F����L%���U���*���`��+�W*ޔ������K���)i��L�6H����<=�s�Cci���r۲����_�z�>.�8�k��ٷ%����Z�݌��#�U��l^�J��eȗ�ɸ�.,�U��7?v��V04���F�)m�bi$ο�>)>����2"�Rx����U�m�/��(D-�j�C%
ۏ��G��ӫ�0�v�^����qiwkx�lo�/��g��rhu��$��__-@��4o�ٵt3�+�ӷ�Kaa��p0�3���S`��I�%Mʬ�~w���,FR����~�_�)%W�v�MO�EcN��jbb�xl���a���V�d�|E}O��=�Vl�lC�Jet�V�Pȉ�v�i�knO�[�F��y��%|�(���:W(J�/W��"ȠF��뚛W�^�rJ�H[ۖ�cŃâU%I�LFDVBH0Sݫ��6UV�E~D��"_E�*u����@��8�~Ǉ�E�̋v��J�|_Gn�Y@���T�+>��v�R�'�Ê�F�#"�ח�׫��wn/*�y��u�ۚ��YV�JJ�ȥ(K&F���"ҫN�0uv�Yr�[��8=��[��� t��ho�����O'��r�ܬ챻���:2!ņ��~K�E������b�e�
�m՝;Vu������j�r��;=N�S����;=N�V���%oI[�V���%oI ��9C^�/V�.��
vzې���՗۳��&��>�wD�1�c&�_,�_;;��64q�<�U�4�/%��}���!���v�9ȳZ��<��P��z��ǖ:n�&SSa[쵃��Tk�ʢo�^������M��U�	�i��I�����;�z��<G"�_��͆����m4��/g	�,�ۯ�K˳�����e��(��_5�]K/��.\T�n߈���p��ۓd��6ܪ�M����*�Ȇ�ʥ�
�˹M�k�i\jӴ����GT䱟���Y�b7p�R-*}4�	��������K�£xu`m��>�.Eo�"�l���g��v�n`�X��|����5h�	5�l�E%���&�6!�Ob�.���������_t��6,�j�y]!:ڕH����D�	�������?�F��dJ�}�Q�q笞E,������Ѳ)6}��_'Û�_�ګ֒e�l�5<^�������wvF��;�]N����T��4R�n�I��R�\H���C�p:�W��$A�u�~#{�le������[��j�%VkzjeoML���v#)%l��V�ߨ�mu�j���jP��R���d��G�u�k�C���)��ht��]��6ͯ�p���S.}�eK'!��u���ú[t{8�Eq\L�j)^��2��b�;�����w�ǩg0mk�e ^?��rwr�Ib¿�FB�3��
��;v�l
t]������{���/F�Nv������I��t�$�"j7n��q"�&�۲ʥ,M:�#Yw��_D~)%�;u/Q�@����ɯq�gWg�߶�d�W+��1'��3�P6���c5��̟���D%G�7+�!VrU�vv;r�)j����a�i6��C��[N��H�1��LC?'�����2lG%�λ�k��?,�Cl�V��/���\�պco��ױ���R�O��I�ݍ�p�x�D*C�N���Sr��`�xdv�/��7e�P4v�U�Q)�%�����,�7;ɟ$I\�i�ҳ��WqƒԃI_O�O;��3��Ӥ�6	!IЮ�*���-�Ƨ_����<0����̅r���P�d��*߷��n�j{?4=�c�֙!I�;�
D����ҕ�+��M�0/å�U/,܁��ï��M�ܬI�%,�B��n
���U$E��1���v�n��o_5�1�=-,�7_c�,��߁�*�c��#�6B�bੵ����j�D���(\��4�ܰo�Ϝ�=c���vk�M�BS�?�d)>�/
��Z��kp����1��VE�����$o��$�_��i�{��h��<������wd6&3J��~6E���sf��o�y
�����ݹm�w4�:V+��=~L�u�ջ�'V����N�[r�ڴ��1}TI[׾?��S����;!N�S���;!N�V��[�V��[�V��[�V��[�b�o�����w�/M��Ȼr�.X4y5sv�@��1�	=ۋN����u�.7lh�ȭC{!3���fU̸�ƪaRE��2�F������L2�wc8�R�Uu��|,���Z_�d�\�8�b{#%�h���(V»ʠd��3���@�[k�7��	4���3�.��v���c}ܱ�&悾��8�9毸�I��M�?l�ݕ��V�V���*�j�ٚA�g�ihp���ݦYv^����A�ҍ��rU�%X��D�H�y�c�����(�ɵ5+t~[�����r1{	C~��/c/�E�r5�̰�ɲ5�6~��=)yJ
N�B�.V����"?�X������@���V��켡��D$�<+��Kѫv�Q�l�X��\�]*m6M��хt�^����_t��6,�j�ys�F�1����gGVU_N���ݾ6�^�7��Y��sͣ�(K	e�����@��RI�a>��'����b$8��gl��d��sQ��=��-�$t;���뎎���Ҩ9;=�Ea�=v�C���}UǏ���f�F���������D��|�8��W+���[;~�)��b��;�����\�[����<����\�ď��i��b���ܑ�?�������/��=��c��I}�?�$T�uO�G�Ҷ����,��QN�S����Y����V�!�>KS*8�WQS�Ys�>��+{��2��'Y�G���t~ۗ�¶z̊�}��xg{Z+ˮrhی	��&��O'�����W�ѻ�2��⍖q���ɨ���]����������U��	N�}�In_e�ɫ�?����i�Z���'��om~.��M��G��{n��R��l2V\��r��e��'�/_��I����K����ہ���͗]�'� �h���vFm-7&曋���q5��w�'��[���b�#{[��6�.��V���P;dW(m��HF���~#���cϠ�`��\��+�ߖ޼VP�w�z�>��^Eg�����p¬dX���{�����$,W'�J���"�9H�&Å^���%�}XL��zĹaJU�5;뷫�6�>ey��]�=��]�_r6�r[sռ�v��i$,
=�U�����vw+L~�c����wh���X2��;��:��9�Y4+/@v������r)���\��1��9���/
��o�iGc�Sv���
��9�ZȧI�T�D~�/���"ut�vR7��g8������|���V!f�vf������yJ�U��_V�fn.H-9\��K�@�	��K%gg
́�9VJX���h֭��ǆ'��ۊHW���a8�X�?ʥ)�>�P��ߵGU	�~��>�7n����mգ!m�X2 �����6�$�Ҝ�rǋݗ�d)�
t�t�:U:vB�*�;![Ⱦ��:�E�����/��η�}o>r�e!X�V�狹\Yv�b��$��`��nBnn����*�K��!4# \��<���	=���{��>z��OA���&��Q	���Rb�$؎;�(��o��]_�Ɓ����׍��C|��*�7n,p����X�+{�jxu�n!#���7[�[\����q��"��I����v��J��i.�E�o��k��*��n��/*`c���M�\�NKQ{?5�qz����
���W�\�.#1�5����P�������W�FH�V9��k{��b^䉱��wD���X�?$�'^&O�a�@���W��J��U������2�-�(,\_KS �E��T���WS�A�p�;Y��X����.������V��$_�5|�vs��뫹۝��2�l1?׭h����_uv����٥�Z�	�g�ri:�


�;T*'#J�ƿ�de�'��˨ݗя^q6��1�y蜽[Xq�/q/�6
Y��_�˴��x�?w�o���ʌ��[8���Td�v)�G�\tz��Ta�u���7�JK�~$�ݜ@x�,��=��NC��Ȭ��q�l?��qOaO�kk5-mf���R�>�aߩ-�+�\��q�O}JK�nr?�R���\��A����/P;�Ǐ��ͳ���?����*�����Pm.Gw+�Yޮ!g{k�|��[J�p2EVP��}JVx�{�>��#��Gl�q����[�6��>݅2P���*}�˔���?�;x��j�e� �s.���;�j�L���g�qd>�qa	�̲6��_F:���ƺ��%7�/!j���y18�5�WZ�y�o�j��[�;��;y��F.˃�r����i�z��,���2����O������۟�ȭ�h*���Y�il+p�N�؍�.Wn��˹萣d�/�V���W#��!m�c dZL_g�����J�Yj>���'��d��*�R���r���R�ee��c����O@�h�ʡ�,���=m:�+-�\���wZ�7���q]S�lv|6{Oʻ\˃�
6Rݳ�o�H2�4ă^�y�k4���D����ʙ)�eʹv�kv���R�Oܔ��wD^6^�,���͝�p���q_(j�e%	�H�n1�����JZODA��i����q�ݵ�۳�S�\��+���$/�/�e�ȹBI�y��sIД�)n���.=�59	%W��kն�D�%	6�_�J����d\�t) ����ȷ��#��\��U ���]�Īa"�ѷ��!��۫���w�D�r{5�?V�7����q%P,p4��"�:m)g�Myyg8�K���e�cr��j�Cc0)��0���)~�Nrn�%X��k���Q�&v�7s��?�1��LJE�a��S�i-�0���4cۗ���JRn˖j�B�_�q}�w)T�V/�ڸ��Y)H��ldCV�ܙ�S���r'mȝ:U:t�t�T�ҩӥS�J�N�N�*�:U:t�t�T�ҩӥS�J�N�b��ӳ��c>�n�jn����'�������5\6�:v)U��%�"��'qF8c�����U��iu	�c�!~p��-۰��rI��$	I�4�&t����P�_��Ҍ��¤�����V�l��-޽pj��ڹo���ͽ�I68�V;�,��V�]�+
(��ʾʫw&��79{O�^f�F^�G�Ȟ�e���MY��I���h�_20����g�k,��ؼ��Ɠ��mUU��n.�� �Q��v11��Ww$\�喵�g�	�J���6�0|��ƾ�VY��röR����+8VOV��f�w ��PR���iZ�b?%�#c���y[]>�Y����W�����>!(H;����#V&�
�i�/%��I�w7�?!�:�Q�.��,��������՗N����J%���Z�	�lND%�:��=�����i+������J�j�͢7��! n!<߆\^�U�'��7ؼ���wm��"����wZ�p4ʌ����z�?���!��M;�-��RF��:W�;l�2��c%���vu?E3k��C�ڏ�H�Wa�J�9[�{A��hyoE�[Y�|��6�Q��*;J�;i��e{�\������698vw�A��a��LS;�ӳ�Ȅ���夌_*�
��)�h쥱�影�&��C��ڌ������(ld:vv���p�_�r?��{�r��6?%$Z�6��{#w�AIkw����Yi���u/��_F�g<�1�4E�&���d$g��]/�0:.:�q�U�c��Sd��"R➯�H��rj��
���MN�v��6#��~W��&�$Cs��g�^vx���-+n/���"۬J�[Ɩܲ�J3V۹ñ��5�-��w+��;l.$X��+�������r��X�%B���`m-�-D�g��`���t�+#�!a�k��V����e�e���xk{�V��l��n����eXH7(J~�E?;����;�t6�G �c3��)>���J쉧`�ITIH`�n���ݍ��&��N���k�|
�j���ϐ��"XJ�������4�i�"���휨�N�sC"^�R��l���R/`�3�w��^N��\�#�)4?gg�FV�&wwӓ6W>�6�&i}Z4e�1��N(���rľ�=��}>�Io���vv����ϲM��g�t�T�oeN����e��&�e���j�~��)�j6��������ճ�
ո�c���r��m�W�V�:�,��с"iIڹ��$���6rV�P�n�3�rX11x�}�ˇQ��j��@��#b��	5��g$RC�I�l��or#��{0�鴳�]�:�l�v���z݄��c*��PQ��nXtCz��T�lD�!������́"H�ݛ���-]y~VӋQ��HU���U;/��7���?*G�H���#�~T�ʑ�R?*G�H���#�~T�ʑ�R۞��-����'Ȼ��e�X䩲�V�����FD�_o?7�O�W�0g@���gb����	j^�ըN}d��w$ћ�kld$�1��;�N��~�j��W�[)�9�Ȯ/�f��^첮<|X��8��D^����o��L��B��.L7Q����F���(�{�e�Rm�&����_r;ui5dO��h� o�\c��aMҁ�װ/H��[�濶���߁܍�"�r�`iF�H��ctK3�5a�V�NuW��pzɾ��ȷk|Y��򵦄�J�9%�(n�7>|U�0�~*&�d߯����I6N�e��<�ffm���T�ݰ�k,��F�!ʲ�m��F�g'�ғ����F��$WP*';P8v;|����;{󤰤�m��`�˥�޼��QN�D��4�VkW``mFD��������`D��D��h��u��2�m��ko0:! p��/��������}Ŭ�9��a��D���%,۔)7d)f�"òP���XiSd[�X��%�����v��ŋ�j�4����&αc� �P6=����oM�[��[+|^P���6���l���G&w_��`qer8r��ݎ�Ce"��J���m�۽υr�,!_piݔ�%#Sr���!�Yr�:V\�����[6�;���K��]�N��P�-�w%��䵶�+n����=YKg!�r�9C�-�2��~#�ɳ���U��ܻ����K%@���)���4';V�NsQ���h���uғa�F\iR_/V�vU�yt���vI^�K~!g"�����iFb�zZ�R}���~M���?&��a�	?�*�?��`h�f�b�-Moѭ�P!\Qzm�K�O�m��wi��}/�����e_�c��û�bi��Y����qz➭ʜQ;�����d�[�|�BD�����e�~W�:��s�[��#��&�H���������#%�[rm\E��,���ud=��YgC��õ-�{Ѷ��V������t|�X�J[��f"�jM{�P�o�5�����)?%�R�r�2�
��f�,�����K�.>�{W�M��M��޼���<u�v�U���ȿgȲț+�-��C�.��)<���p�����%,��.M7g��%'����Q����?�m޲��:�\4�*������@��[e"l�Y*�y
�7;�c�ό�n�p��Uw}�����z�� qrzufA��qK7a7aR��HȽc�^��vUj呏��޾�-nM��m�W)BR��S�u l"`�	=�_�3g�&�\���m�W6�_ ��V�헋S�,�瑑/!o�vB6���g<�Y蒻8���z1 t[`�R�yx���O[�����$�U��߶<�T�{�����`�H2�V~.+��TnE6�9er��k��9�T{2*�v�$�J��[n�m˜7����#�~T�ʑ�R?*E�Q|_�E�Q|_@�B�TU�^�7"|6hV}Zo�N"˃���nn\A}`Ȯ�v��`��]���d�,��K���"E/	U.�	�5҉.K�s�w%����.M��h���>e��%�����ݖK���Z!5z�\��Se��=&�V��n�vI�Y�,kQ8tRf�I�ך�z���M�����ܤ�eP��8h��a��"Ý���s}ݓ�}���IN��@���'�n�p�35�\p����\#e��8��K�}}��Y���������y��I��s�.R~�+������α����V����'�%����!���od�˿����丬6����Z�!��\Y��a}�팍l��"����n�tu����ϳ�׻k�WJO���E_��V��M��"Y�c������U��y�^U.�S�Q/(�/Vx�_Ϟ���?bp�F_�		��Y�&��'�*J��.ѵ��'�<�K�ã�o�=a.:�@�����������j����U2����w;��H[8�����2�oY��c�:}�c��rv�n#�w8Y��{�4��Q�-��H�����ҫ��>�Wa��A�=ͮ�s�j!����L���9����gZ�p2E���P�|S���u��kQ�-��k10�E��C�Y�P+Q�c���2R6^���[��lw�����6Ƴ��[%-�wQ-��Mk���_e�����|1����N�ʳ[�T�P��b�A���"d,G:b�A��6[-{l~�;C3��e�ޜ�j�3_'�W�s ga�,h��U9U���@��c��v��j����Z�G�"u�{�uh��Z��]�P�[��	f��dm������2殾��m��3n��~�^������@�`d��ͥ�}�v_�ͻf��mb�$YI)�	W�E��(��9��K��(Gd"!'o�%Z*�Rir���u��"��7�ON�P1I~!�g�g���BG�y2-}F��c�S����]��=���W%�Wu&��I�R��'�.���)H�#�]�)��JU����'Ca,rی��(��}�q�%�ϗ��n��w|���+���O�����m�}��;���������F�d,���6��L�ǥ7�$�`��RN�!"�o�1vx�H��^eWȹ<��2�����l�B�V����se��\$%k���U��]����nR���Ei�a��]s���OVۻX��2��j΁,���ȳF������݁�S�;7:�g�׳��&����wE:�_%m8���-���g�������ɵ��O�d��ڔ"�T+'��nqS�,��n���Jۑk�X�W�eW~��o�ZqK�t0Z�ݽ]6E}�&��,���"s�85�&S��wW"�ϭ��£8l�r��/Ir��#�MZu�3_��:�'���nYߑܖ-��!�7��o�����?�|��������N/�8�����N/�:~T��B�g
�p�8pg������pӡ�����Xl�K�7VE=|cr^B����r츍�sQ/h��
\>e�����a���7;W�]��q��a�,�,�qg���r��s\XQ���/������ݤK�N�yEV���pU�K�yߥݸܤ͹v����Dg:08p���M�Eg�{Bg�l�Y�܍���p�����ю����f���=z�MV
Aߓl�+=4�,��c��f�hW�XQB�Q�go*ۇ�r��J]�9C_SN���F���r���4����=d��b)Y��m���|���ܵ���En���n`��*���
O_,����ۂ���$nûْ�`��h��!. d�`y�U�~lʵV���J����g���h�II��Mō}�a
5�挰�	��Լ�񱐑��9�њ&��O		,���RX��X���n\���+����U=�����M�����o���j"��*�ݬǲ��<�n�V����-��1�b�M�����8��t��H������myz}8��s���#�2�+#[侢���Eed� ����n�t�5���s��[�~���uSS����1��m{�����%���+Y��DS���edv��I�)S��ʌ���8
}���(8�f�%�Qݬ����P;l�/�wk��P��*��g�V�*����<��H�e�qy��*
�M��jt����h��5�|k�����94o����e�z��K$�YyL�S(Y嬻�9CJR������⍔$����A��..��L�,�/�:��e�k����������'�d`n�!%�d[����z�Z�l�ɹN��܄�G�Ѷ�xN-�Ka[+޵�ߒҰ�IQ:��Zܫ��֗�
n�+c���g��v�rP=�����x*���=&�!�L�p�dZ$�[��^H�wa����P��,繑&�$��bO�����ݬ�IJO�l���mIZ�O�ܡ"m�wt��
KЇ���-ά���tr|7�9+���+i؋����VuW���}�6�/?��ّO���{Ve��*��ݧI�-δ	cvΦ��s�o�ox�{�)#B��V��Y/��'
z.^v��}��
��b,{���H�m$�P�����e�Gӆc�m��������o4�e��A�����ȣ�ϑTeZ���ߓV�������ˆ���X����V5jX��q�@9Q�\�	__-��a~�[\0��v%`�ȵ׸��K�׬%�fD�6��rU�
�a!}�����I�.��&���2��n�_i��\�5g��/ɟvA۸���dU�jˬʵb�E���|�g����s쵏w=8WXVC+'i����*	�N��HX+m�{�X�P+�P�%~�����_FD��&�?��?��"�!�|_q|	�p'm��:�v�	�p'�B��+�Cl��46��*rJ���+!@�!X���'m�ѐh1ˉK^���@������ǃ^ݰrI�)��(,X�dg��n�_z�T�g<v�L�g�5�sFY�0�E���t���i3Xn��`�hRdu���H��/~��Z,p\�Ȭbs����*,wW�}�a�'ZD�ɡYؾ�?T��3Ś����� h�E!�/��4~��qX��}^;M�k �X���>��Y��d\k�0|��!V��o����Ɖ��V1cj{�<5>�iKr�e�W�Gԫ�;��_MX��I�ڋ���$�e�JC��q2���?���Yړӻ2��D�Ək�P��tC�v�W�#t��E&������`X~rK��N��3�j5z���B���}�J%R�yFiz��j�|��FU��3"Y��q�&�De��u�����&�D�$�?�����q�M�&UIa"���	�_���ܽv��/EwSL��j2_{�H�O�b��EG+��P$n/M��Ǥ����<�|����z8�s�� ��R�m�^^���5/[�q�
����Ȭ�������`����OH���uq��Pb�s�������j��S(y�R+#�5�/Z��5FGwi�m�2���Wt1��z{Y/�8Ҷ��+���-�!ej��Vk�^������Pd�sZ�J�iZ��"��")q���:ϱ����Z�KpT�o����^,�[#򀣄��\+�ZQ�~J�q��Kɡ�W��+#����[�����e�BH���K�df�i=X�K�R���P,�Z�l�?��0,�?��}�B��9#.5|���&��T��Sm����:9)������w���0�̾��S����OOS,�E�	c���A9�����ݓ�AUՒ���)�m�c��������ݦ���ܻn~�-�9CK�+����P�T6�Y�D62����KY�W���e�k����)�d��Ff����*��ɱ{�m���i�19k��d���:)�܎7wvG�EzY(j�鸬�~y-)yϕ�۱{�!I�04{b{5=�V����ۉF��	�Ue�JRv�]��4�o�l���8�,}ކ.E!�V�-Y
E��a���qq��_��#D��_���v��;k0�/n�~^����I�kw*�%M�ٱn+��g>�v��$�����l������#��?c
�R��f�%nYjU|�_g=\�;������g��իm���[��@�2+�/�&�m����������I٬��I~{�>��j�*�iH����U|�q��F�p�Z��
���vɤ�{~o��&�g��8�_.�U2>���d�Ѵ�I�&��kȩ�8dLv	�9BRȔ)��l*2/���U/r�nK)2��H�y�&SdL]���UF�w�U=���"�"���t�
�p���|�n�g��'rdQ�ϫr��^X�\�W�`Q���"�iI�M�BB����"r�^)d���c����6�ٓ4cZ���l1��s�,ud�{���n<^�%���{)ݗ~Ό��*㤻����y��݂��/gW̼�?�
��O		_����AI��̪ZvP5������K����5��m}�,��U.l|�9�*:�%,��dREbQ�B��YfK�Ʒ�c[��r�dh������I����7K6ݚ7�3ƭ����ݗߑI����(���ν�%&��&���I����w���~V[�·�YW�,_'v�#gi���Q�m��F&��ĲOa�����'#K��Y�_K
ȋ�y��%�h��6
���˷���}��UN�볝�vr�g�]j��c0r5aT
�}��@�聤��7Y4�K����_��p$�9=d��0Q8�}yd�����Y���(e��4V%j-�K�s�yzUK8�[�[�"�T�ψ�d(��59N�������#��.|{���G��|V�g>��@y�@��=/B�����%����s�����ƕ�ʔ1%��ĭ�A��j�%���V� �b�O�]��JUqZ��zվK�d�=2C���m����4���Q��-M+S���{���+��[�)*F��5����+;���c-$[r�O�K�@��Q|G����׋�Pܷ���"��
��e�6KY��?g)gQ�ȝ��]����]�_������g_�>Y�����I��nɲ2P�V��V��}>E��V)�,^';&� ZU��xU��o�=�>*LF�RȬg�+6�?�I[y^�|?�����x��6�5i����~�n|�~���$������a>X�,��O��4��Pݼq���Z�*��X�5�~�VަB��Yn!��2�#-@��b�U�@�ׂ\�`����M!q<����u�d��ҷm4�6�V�A���BH;j�c?�r'_gX�����m������v��'i�*�m���U�|��h���׻C�rx�DNRږU��J��G�߁���\�j��G;g�`|o`��3���a�dfY�dUX��}��6������Vv�[��{J�f��'X���⍦V���[�,ٷ<�k��Ձ��դ������@�A�wq�h�f�J���M�K|^��,�ΕN��gYy3Q,��d� �"�aڑ��xPLrj����,^�c�ŕҌ�ABE�
T�M���ʧg,rg��i�aQx�-�rl���߷ �l���KcN�P$�,2�w�,�ȗ�,�7k��'�ǟ�����������5�B�w̾~j�Z(��ǯq��>A�Ȳ��es�k6��v!J�nY?������_�[�ݐlm�V#�����!P�����W�I��e���*���|Cq46�N����vBȫ �K�ص���>D�7���:�&G���2(�,��#��^L��ݠdUݖ;$��;>��ȱJ�kf}��:4�6z8e^{x�a+�㌗���x�106�����ɥ讘J��4�U�Y����x�������!o�ܤ�2.�D�eTC#����nk����q_/j��:#t_�̿3��\�5�f����n��,��Ыqv2Y�E�8��s�I�p�ga��MI[�d\<�p*tjA�шȍ��j�c�Wc
�IW��%Xn©9Ӭ�qz��n�k~L�\!*��_��m�+]��R{�<�)7kp�2xˉ4M�?��+�jx�{-ƃ��!�����i#{Y�[��K�:��mƳ۴��R��$g��v�M�HRW�^(9Uؘ���r0cx�.�]_q���n��Uz�^_5���g}[��ѽvwh�}[�j՞{�44h����&���g��Y�������_"�ݹRF��������dO��ۻ@�K0p#bby��Ú6ϲA�z59x���ʶ�kYZ�F���(/mcM��m-�]�����I�Z�Y�����vR�֥6RP�I,�/唥�i�\�ky������L��k5,F�+���~YJ^&;l$�6����ַ���{c��r�Q�Ov���[5��f�gS�r��KY!�=͗�)��G��j}A�����W�=��Wn\9��V�[��i#c��wi�,��=N�Gem�ۖ�H;J�f���Kp�?^M� �q;�m�*F�c(Whu�ԇɭ�X��$�" ����'.�U|���]0�@�O����ўd����lC����썿��
B�����ؼ��a�"Ҭg����l���҆����ݞnQ���݌7R�ß��^�_̛?ϛ82)?$�3�2���M�'���D)��������|e3��x���>̋
�'gf�B�)���E�Y�D���jr5n;���ܬ�-��l�3rO���˯�ֱ�b�J�n�����(�ǳ[!I�.�#S�J�I�>TmfP��T�~�?a!6�Z�cv1y<�e������_�\]i�B�MqV
]��I��\�ݶز�m���o��콶O#V*��ܕϻ(E6WӬn2���YL���`UYѿ�
��K���t�[^&H��T��m�6^ �g��Q�؄Ӆ�i���S��9.�{U�DB3���/�c�~�E�'�ȁ�W�����������R�/�FA���n�*ğKc@��Β!'��F��Y�FRU����җX�̷[����%j�J��#*�ߢ��z ��V��f��œ���v�{*��@䬸�������AW٥Q���u��~I@��on[��>�"���ܭb���4k������jx����g�ń*
�2��c	��}���Zݟd^O�@��r�o�����e	3!���׈lnX�L~�����ʳ[�l��,F�B�_����/�g}�E~�����3rLܓ7e�)b�^�W�l��Q�g�����X�X�lP�;�E~ܚ}�w�z�^�Iߒk�$W�I��"��{�Ƽ��^��I�Z���wf>�5�	zK��c5�W�.���玭Y���L�}_�'�]��Ѱ8a3*���K7$KLq�"p"pxe]��2UgɁ�M���7�~�~��~ᗄ��a�z�0�3�$Z�x)?�mQ�5T���o��Un%ז��q_Ł��
*��w�h��ݏ��Ye\���������cM����7z��Ӓ&�R�BG�1�K#-��r#���`���4g�,4Zݱ��gc�����dB�Tcz�ߌ��S��j���B
_\����P麙M�����ju���۹@�q[c��"���K_�gnW�m�ՖW�H�I����Q�k7��y�Q�^��e���o���T�Wh�}[�j՞{�41�K˹��,�W����ș��n�Rn�FW��%�{��-{
�c�Mȶ��)����nie�<��R����:�K/��)[�Td��B��d����n�-���R�廟�����q�W*eO��x,W���k\��ޚ�Q���)-�Ij����4�e@�Ǽ
��~���w��K�{\S��{ �}*�ۢ�bټ�C���V�%��GQ���)-J�x5�K�H���=��\�T�WaJ�u�5�+��ӳ��en�d�~�nG�)_��2���ä��GM��֢��v� ��D�q ����n=
�g�w��nwe���K�\�i;rZ�gg"�%�z4o-a����㬊��E�:H%��8��y�'��̳�K9�,*ܫ���r�FvRJ��3D)���m}�۔*E�2v��W���{��ۿ�v��d� �z��f�qAY�D���cwcdЬ��?'*?��-�*���ɩ���NU�^ƞ�����ق���"׶�g�6�������ۓK���H;��f!���]t[r$�4�	�Z�JN(/�:����f�h�K}�B�vA,���6Yd{�_!�#u�
��*'e�%q;<�U�k~�z�Ic��X�/�O�0HK���^�x`��T}Չ�W4^�η�����V�����5�'��aA$��w^V�\�<��f��C�H�VY}N�N�����\���
K��M���HVu-��unƇ�V�عT*�����a#�vv�TN��FD��%|��ډ��D�aWkv�57�rp���~���_��q������IP5Ġ��$o���M�e����^OF#��F�~�Z�5��up��e�z݆_d�������^__M��)`K,<�/�:T��:P�6r7欑@�ၧdZ䳗�XNM��~'��ׄ�J��c%�1�vh���&�RH�#,�>��Fȴ�XH��g����
��)�7-o$7��e���[���#_�!��	����4�>���Rfܲ��2+�eWy3�ܵ��ia������H����������ȟ�k�dW�I��wm��v]~r�8n^K�cnΎ���xeR�x2��fzY^��D�$Rj2��G������vȘH���1����2f9v)r��r�7��y�a�_wE��͌mc����&�s\X�*��G�����W�Y�N�J�W�?4���+�T�c4K����?걮):�ʨ�'�H���H��f����ȾE澷�X�5��a��0�n�Y�۔&/^����m��^��I*�Y�����,q¬tvج*�.�᳍�n\m���5��|1�)�9�����J�e(�O&o�����79*U�J���I�[��Mx��M�*�z9[��K;m��	c[�1{L�^�����k��o:��=��O'�����0�������z^���9z3�W=..9��ϟ;��UN�Ev��ջv�Yᗻ�C6e�K�y�lɬ�AF��s���g&�II_g"������ϭ��ʥQ���mbU!S�qu����P�ҫ)#�P��*>���H|i+'���M�R�W
T��ۤ~�H�H�)C���q�ͯ/Q��vͭs�{ �|{�����ĭ���f��C�zh;X6��ë��{�����8�ë��R�=��[���R��� ��K��T�s��ҳ�N�����k�~�;Q!m(u����|H;H�;[�m��JU�g���{:�˱��i[ϔv����*U��l�l� �%�N�cݻ�k��b3�4�
��x�[i����ц_��Z,b`�d٩ ��Do��<�/�pʣ.���² �_w��i����)5ʒ�U��/*��Y���7�*L�H��p]����7����ݸ���m��rI��X�"�ɝ�h݉���JT������۰��X<�<����6"�*�SV��XyדqV��6Zu�-�iX��x�8�rU��/���LN��/��=���w�Y���-[u�8_g添�픡5�t���;��A�xun1�aʏ���I+m����k�|���͗�p�
�
�
��
&hB���,�w{i2��� ��G'���n���rKlkw_
NI��t{ `���Ϣ/�[@���.^Q�*%')�$�9-Z��6���G�wͳL��:�K�:M���,5����λ�R}x-|���l ��Y�4�>�J5���~'M�j/_�ݬaՁ���V���V�v�W�%����VVMVˁ��*�
��E.�Bi@�CdQ�w+���$ߔ	>|*'^A�\�����mF.,:Us�}����vJ�S������m�d�2'����
ϷG�pg[��X��a|l"61&�Clv;u�V}}bOr�	"�&�&��'�K��Ul%�|�<�ξ	��_��w'�lw<ө*�U�f�����$������wp$Sז_�^߰��#�UHҳ�٫k__6�E\�bUH׍gĲ>��vt{r0�`�ߑQ�if���b����{������{��-z��ػ,vtx�Upl���E�~<�ט�8DN�(ۍ(G��*�`F����D�^���yu~�4j�q�6&�1z�:��u/q/�3�w���s�a�N8�������e��6M�'�w���p�ї�v
O�
M	qI֏�j��ga	'��ȓI[=N|+�r���G�_q@��T��"/!�0+RS%�����)p�#��\�&�G��8��O�����d��U�6��]�Xݍ�qZȍ�a��Dl�1�Us�%Y(R�2��u�Q��r��؅3	���m�b����B�����\�\2��y��D"�Fw���~�67���2!�ɴ���hpdQ�7+����:7�^�Y}�\\\s�F���UN�Ev��ջv�Y�����5���}|� y��D��>�c�I�e��<�M��6O�����co���0�����o�}���b�*�/8��b�d��[���ݓ���o�[�T�G!áe��P)r;�\x���g<w���0�usR�a}�)�1H�����צ���H�g��o1Hݜxv��� �~�X�/Ƒި�����<<o���:w9���b�K[���}�X?G���I[�[s��U�VK)��C�P���C��H�+���5�qZ��:쬬�duj=��$:◊B����>���܏��k��[y��� 1Z���Lߊ�s��1�Y��2�k�R^]F�<���ݣ4��������,~�����%]dPR��_��0\80��pW)��'����H9-�Ȅ��N���[q�^�BP܂��U/M��<���-M�MM�s�������	ٟ	���%p�19]5�>w,�7�J��ke<�:�i ��$)6�B���l"�$��fmyf|�X�� �4�1�4���d�?��Q�烒����R��ԃg���ב����Eܮ��c[׹z$,��c�!��S�H{H*����m��Z��m��nEʋ��*�7:�����݆����s��v���h˯+��{:n}��H����^_E��r�9��ن��'�l�*�W�wg@Ҳ��ߍ�!g�|�7P��ԖM��c���c%�܏��g9Cw�*c��=���)X�J�ȗB�l�v���YjY�c ����V7c%��C`�6V���{>�8U%cQ�ͫ���J��Y���in�cey�/?]F��,�;U���ո�~X~J]��>(jܤ=yE@�����z��*�)x,	�� �v\Z�����'�[����2Z�2�����UV��'"+!`ٹ[���vx�%�d�$63��M)io�y8d.̎(��5�	<�|���B���@��ξ�g_�������i6��܋�5��ia��ë��w��奣nUknEWnYv�b�S�"i�BA�i������+;r�I[��CW�#6��슎����^�&��_8��8�Fj��e�	ܬZ�-+䚎}#^ŷ��nUk>O9�g��L׋�ȷ sD�lo����Y���X���quD�WD�^�H~z(㵏�5��^��=ToL�W6��/u��c��O_609��9��[�.J�$�J�&E��fl?��D愰����hL>i.<���J���^�5a3Q�i.c�a������,ȶ�1�^l)ۉY*/m��}�kv;�B��Q9�/&�;~���'�G�'��Y�'�����\76q��%���TV4�n,�D��U	E�k�X`b2~I6/SeU[rU��[�	'���R������4����-�uoΖB�3s;����(��+;�sF����9�L�r�Uh�^�\6�v��T�Wh�}[�j՞�4�)#3FF]��/ik5&D*ˋc�	�*�k�XYȭy��,����܁�דG�]�(����g���ʶ^��S�O�j�\x<W��g�P=X����8�)���w��������/��A����;�?��g��x���=~?��m�tq��x1-b�c��x2����S��~���\�俦���;���x��s����Ȭ�[�u����4�>�l�ժqY����vK��?vƳ���r�9Y�����YO��2�{����2+#�Yx~WgQ��m�<�KaO�j#�iC���Y�]/F3S���e��6[��������IG<^/K������2����.��F�����c�p8����I��l�m��N�V��J������>3>7e픫4�f���F����6Y
���ȵ�o�曋�;rȔ���a��r��啉6�8�f�L+/)D�{��V�+.�%r���&�m�\Sw����j��nP��e�&��;٦��!���bB��xdЛu���X�'+�#i�r߉��[9Vv�Lo�A`�s04Y�k:�78Vv7�q�����dX���+I����Cީ�	c�&��/��i\a�@ݯ��E�{CFG����ɨ�Bet���k��X���츫M�m�e)�u,ijw�ya{����V!,���Kܣe��X����O^'��s��K7��	"R��\�z��9��D,]���|^h���$\��|���e��m��f�f��O���Z�}	5�Z��	K���X�d=5Z�c�kw%��� �7��¡��'5�7R{�5[��5�)CW��&���t��eˊ/a�[�d���d�!\���v�yח��b�J�v)n�[���F��D�w���S'�H9�R{��srk��k�����
�խ��b�Q/CE�I*����brU�l��_,�oʱ5���Īk3w�ܞM�Փ�dQ7(�
�2j���wb[�]�MzI�ɥ�0q�����ͻ�ϋ?7&}�n�8�XV��v���۹וfՓ]�K%�03vX߫Մg�d@�!0ITk���|kV5Ɂ��U�>MVU�k?��N���_���_���J�qJ$
'�X�z\�]a�.���r��4W�o�����D�QN���:�=$��Oc�&Y�Y�_��TL��c�W�>
M	G��RhH�o>��9�c�F^�XL˫Q�eຮ�����W���D�&Ԛj����'��*Y�.�Y�H�4�;r((��J!϶Ύ�d��O��~��cE��쉁�J��PH){�t!/D��$X8��|�蚫hڨ#K3^?��K7$\�*�~�����D$�L��-���?��T
[M�_J�����]ȳ��HZ�iC���ƖN�%}&h�(�����XR��8j渜�[���(��_/;��gj�ld�Ý%#��Z7�������3c��`�ʰ#s�Ul)1�g���|��g���cҕO_J(Xr����Z2?(I��6Jܬjy+˕;��������X�ĕ�ϹJ[pܷ�;ia���ی����ȵi����.������䒴��X:��>���M��V#$���p�d������o��"�*���C~��#0m�:T��Ub�>�a�M�����«��������JA���W�Sr8���,�~|�,ϔ%[y�͔��R�re{k{JƲU�e�J_�m��H��}�����N��]����-i�������E�82&*,wW�W�F��1�P�rx$�'���u�\U�,��"���`I�t�h����)wr�ȯ���G�w/�y����E�Ҭ^��;E�Ռ�����:Hm��5�f���B��۱����v
O%rF�4~`I��=�i�c�gINߍ�3m�ȩ��i#{�����O�c���iP�Gv���6/�����n·Z�ili��/8�nT����u�r7��n�#M��)���˼Q��,d�^H�Ua[�rK3Cu`���sV��>�b�\p��L�YR�.#��&��p���Kg�[�%UR�Z���
�C��Nܑ)r[�Wn]W�l<�\ָ����.7),m����;�9��is���Z�K�VY�7aRd���Ij�����R�[�BY)m���u�Y���I��3�\�qyTB���/I�Y��-��g�,��Γ;�a�ۑo%��{�ML�2K�%�[&�[U��Җ��
��_��Z�s�Я���Q�����;���'[����T��[�nH�a,8�>ʨ��v{���T%�/��qK7sJ|��=�����D���m-.�]�~�RW�$��>s�l.V+-�^���>�(oʩ����B�e�����Y�Ȗ
7.��[>����/�������qy	>A�`�{k���;��s�gg'�'�Z�v\\����89�%�{��+8$�%�c;�,|\�:����Up,'����ʾ��]��ܱ��aW��������/��I���'�_VO����n��V��d�Ϲ��/ϋȤm:/���(�\9��/�N�ׯ�F�7�����g���ٿ滎�\tn?���F޾����,%��c]��2_�q����Ưϱ������Nh�v�����U���Z_p+�Q2�d��K5|&�?���237=+��6��V1/���;)F�gŃ_ׁ���}ǯ�^U�6�X˔o�/6�����Y�'�����i���g����D>¤H�6�u�2,8=e�])4��e�JX?�V���锝��:��q�XK�Fiv�(,��g�둂�F2�����溾%,���X��a������捤�����D�h�qc�
	/uU:��+��v^��U��̲��%#��:,i?�K.��u��_`��׳J㋱�B2�O�s��_F�}���X��Ɏ�[�Hp��M)m4��M�^�~R�D%G;g�m�pӶ{�ݜ���D$�7M#ev2�*���[v1
��ˈ����![��,���K!jd�+��9T�Fҕ��[���~�{o��Q�6�ߴ��r[Ku7;$HZ��al�Gx��{���������>2[o%������)��r��/n�V%)����:��SaZ�wdn6��e7��T��S���sL����������c-ñv�~��$Kx�$~ʔ����n���s�)B���E5�xW��Z���5��|汉�I����_�	u޲����*���������S$.Jn�/���T;�߰�	3KD��,�\�yP�-O���r1��]]�),�2%��,��=�*��*A�wm�ܫ�X��?:�h*�|�Ã%P$*f���e��ܮS��������U���qw�l�WW;@���2���^?�����m�[�e~��k;r��P�����X�~C�7���iT'Y��ۦ��G�{�|�歳[c��(��I��_����<(�U@�	z�f�!�+�@��r!�I�cj�/a�`�4��[dSߌ��������	��aM׿n6�*�p����j,��&����)���"R�|���2���Rl�	6#�77����[�]���K��^��;�f����ΰ4�7%2Aߩ��L�l"�
�m܃kTd�!A�����^�cU̗Q�τǟ�_u,�pgځ��V9m�ſ;���r)�z��=�l$���>�F�$���%���M�1��C�06jv�,8}�y϶�%�K�#W��U�J�M�"۱ݬidV3�T��ȅ��n>�p!"�2������K����o�Ss�����	'��!!Q��8H��UV6�c
����+�{;�^LzVx�ƣ5y��w{w����*�X�j���&��g&��WѕWѱ�RF#l'_&��"Ñ'�����c����IVUۑs���|�%g:���d�_>�^�I~#�F7UX�v5,�I��}}��2�a]�;�������l�%X`�����F|��D¿������]yz�����?�``cn1��G��tN�ϵ�����Fs�D֐4�cl�4Af���}�fl3���b`e�n.�h��q=�
!*��1�gFUWJ7[��"}�q_&�����y���,����az5�~����Ywv
E(\����S����<�a�g�M���ܳ��n>�P�W�ȶ��G�Rʐk1��7[��}��;&��B}��ݸ�ȳ�P�Mv����i.[�d�%|K�?�{���+��Z�Y��֬�X�MF�&U�_���E*�����K��W���ګ���=\�:���'�l�7PP�w�K�l	<�M%J���~��BF�$�{x=��-����[�6�w�Q#���w������:����6�ؤ,��emGk%�R��(|tS���Tx���Y�����E!dV��~<KW?�k�xh4�^�R��R_��az�V��|�;���em��Px�Z����v�Z�K��������x���Q��jճ���8�5O8�Px�j�j>=��v)���|�2=��r�,^��N�Hu�������ڏ��JH�v��NN��(e�d�nv�A�e�/�H�kdiJH��r����Aoӝ��u�n�]��jp%,F<�ח�cÆ��7o����	��B]F2o�j8a3Q���&o8��y��,�My=����Ěۥ��d�)��9CwD����*�m(����WVP���B��w��7~���$T��d$�S@�Prx�U�o�YZ�Z���H��U�P���[v��B���&��ȓP8���2�d呶�X0Q�8	fe�:���q�v�"�&'e�"�l�\�r=��i�V�2��>�}���*�m��w����c(_�ܱYr1�-�rܘ;n~��s%Z$��̌Gm��}_���6�2hɣTw!�K{.�ܙ�jU�;32%����Y]�~U���Yw�x���wR���ϲ�eX��V4�W-����+�o�Pϰ�HQ�hS#�Y����r���o�7n���\Tn_��FFG��X��BC�ea�L�^_�����u�^�f?�/>�jVl������kw���~4	���V_Dl6Mks��H�X��S���]�U�W�Sr���}ܸ�*������z!�q͆Z筌��&��ֳ��+5򔋒�'�J��^�^Y��׬m�k��i@ՖUW�X���{v���O%q�I�iH9����y�Z��F
�'����٢��'��FդU�c�y���K��0%�n���r6�2,���&�H�a�q�f|^Y��g��M&��WݖXΒ1_�F�cg�<�&�m��X?Vݕ�����}K#/��X@��Y�p)(��N�Mkr
��N}�D*O@��$��7z+�$�p6��݂�ƞe�r�˥�U��R0�J��T���&�hϝ��a]�v�9z6��U�3�ca�I,ϯ�_�4%�q�D�����<��^�h�]���gk�9�}�k_|����,���uT��2՜r��"�&�{�W������(��	T�M�Y�U��OÃ犑&������N�D��v�V���cr��_>2���m&����T�/��_�I����d�ݥo��Y
Ҳ�q;y�xVw%�%b��ʜ�3X�¥��C���k��ʬ�2$_ws�n�c���gg'^�ל��mK��U�Ѣ^&6Յ}��
�aoU(�Wh���5o�/������i����zݸ�s�I������JT�qx�_J_��� �%�H��-�hW�Gw[�n�`d�Q:�m6�񿴥nedm��\S�^�K��:���"�P>R܎���[y��h;�N�#���S�q�5sS�Ii"��{e�V;�m�?;�e�?�=6���Q��h�Vä|/C�A�5s���K�!�_��{+��[A���t�x��/J���\��W��S�����3y�xI�.}-f���Y���}��l��L�N)whyKgY�╍e>������]�}�.�[-öqX>ҧ����gfʙ�����v�����B6!m�'�*�_:���Ѿ�Լ��j��yɣpȣ]e��OL�doZ��+�7c.:�RAnɐR���>�t�����gMrF�l����I����a⤑S{%T�x�J�5�J�!&܋�ܫz]�nt	;nF�wce�dD�+;-��#���ا�BF�v�2�9yAdA$_�T؆��9���n��nM,�k��t�$��sD7J�r�P�L���{@�e���n�VKp��k/[Cl�P%_x���Q��7�SMY�FޠX�PWӬ�RV��W���$�e��{0�3:�P=����B�T���j���`f�������TZܫ���١��ҁ��>���5�>���0~���`���'��g�)&�FN��o^�������`I�~�`�ܰI�K���rI�¬�nF,f���]m�����Jȗ��P4U�����[�bO��۰���mS8bk1w�R�%�2~pZ�WP�\6j�BMU���)iD"�i��6J҈|����;.��94��]�(H�"�V�w�n�s욁�)Ն7���MX��g�N�B�w�2�W��c_����3�e���1��0[��$-z��n&_��?'���q*��ry�f�˭�*���gk�_+��eȌ�����y$�6�)k��p5�;r|���ܛcÁ�ۖI[�9]��#YÃ(k��$��(ͽ�͹T����
x��)��O
r���_�R�	y<L�>�Vl|����)ȣ/�W��%\困��T�F�M�������*18WU_�|��Rl~q��0~�iX݌�	*���F�ر�q<p��#9�I������)T�sKsW�U,����ǣ�-yޢ�5��zѣqv��q	_��Ļ��9yxNdV2�,���ecn�&�����={,P�V��7��#Eڸ���,eRj����˺�u��I�dyI��ۉ�����20�,��:��hU�>M��"�w
��#_�ޢB��s��c�b�����H�=|�A�"���z5�����:Iy<o����ȝ])��c��@��1�5eP��zt7"/��Ea��5��4�5u|��]��G�34fZ�͡q�'��ԺuS��Vwp�W���W�@�,n,)-FA]��q͛3Fo<�{�ݎ��{_�ʠ��{���d6PBK"kx�L�gK���i��m�F�Q������;H�d���R��?�sC�A��w�/!�x�S����t>G���Ʈj0~��%����o��J���ax|��o3�׀��r?�� ڔ���xk#�P|S�������������q��B�+%������9�C��N����^#���c�A�Iht1�����x�K[ΎZ�:8�zG{�O��t�^��������� ;|?ǧǤ�7;�s��K7eEk%��ۤ����+�F�F��]�9K{cX�K-�Ɩ��U��f...-c�q���.�ZR/��s�����W��q�sFy\ac��5Ċ�'�#�YM���FJ���zB����l����W�%U�M��"�Ҧ�~i��t��V�r1�!�p�]܍��%v��h�nQ�ؼ*ݽ��l�2���nU��ִ�󰦗�u�N��+\Vz�(�E7�ܛ��J'�!]c�PRld��!r�DۗK�ZʣXw��T`��b���m�a�wl��J1U�q8�T���ȹ���y>�p)7��)� �2��fJ��b�Z������2�E;_�ÎU�{Ac/��o�7n-p��X�M��C	p��I�7���('[�$M��ٴ�~�n7�$��"�ͥ�sdANM�I�-n���Yɲ\�2�?5���ܞ.,X�-Y3-'E�1���c�m��u���P���Q	m��@������U<�~�\V�2;���Q����ȥ��,p�v"?S�o���Ww�*���v{b�4�<�$j��C����:�c[�����Y�D�r&�����$W��ݱ�O�'���	������&ᔻ28cs��,3�F�fҦ��IY�y:���w2��0�+X�ݦݟva%j�P)%���e�c�����{5����M-������?a[�h�RU������rZ����6v廒ܠJ���E7�O�߰��vU<�7Ԫ&�)��NUIFEIF6�W��@��g�IW"2슒��M��4$�f<ц7:�xf�v8`d]X�j>h�qw�1�t@�L��|
�7^q�]\�^`l���UT��	j����h������0Z4yªQAX�׹dX�F��$�]c9ㄵ<��� �]�F�u[ז������׬k,���*���I����Dգ�	��&��*�[w �d�a3*��c��q�EX�8��v�:��+
�w>��3��1��<81/�T��۱8�vO��D�ݲ(܈�I4'$�
͑��'�d@�#p����&��pܥ
lC-%p䬹ժ�~����\I�?���Xu��n[h�X7����ω�KS�z��n��j_�Y�\1�a��֯_�y���_.�/}We�U��^�]�~��W��I�X�K�}�		V&	�������������ۭ�ۖ���o���<�z������T�d�J�����+i���w������[S��2�:�[��=>)�R��,V� ��݊{������|���|[Y�?��z>t�ߩ-��>{��K��������Y��q�s�z����K����6�K��>H���n(t���b�?�Q�)��R�b��-S���qn����Vl���R��mv������%�r��P�w�H�����ݤ�ɼ�ܻq�y�k|�S#`�*v��%d�\�d�!îZ�n6���f�Z�����8��tQ�o�z������.�E���v�<㱄�&��gc��3�>YMߞ|l��DA�-����)����m��IaÃ8�;�^�E��޲/,��ھ`��f^R�ki��9)�Bk"�Z�m��R���F۲Ҕ��G��f>�o��j�r��,��,��a׌��Uݰ�J�]��q
��X߯����y��S�U��C�5n�=�W{@�֡5�5��6�yxVO��z-�{v"UA�Q�����;t��R��x�-�Q'��]HE\ϯ�rh�m"ꍗ�J��B�V�{(D���!&I�����~U��nP9�;�7d�V�(-ZL�zL,g�9fm.}d���3W�c��"p�ں7bd�^�D�I)~3�U�z�X,saױ�ݱ�����,���|����]'�>��zl��=|:��r��v>�r@��QI�����?w�+�ݚE��������^^7<�-v{>�/�܉�܉�_w�'�A�l)ѵ��Ҭ12~���HW����,50����qX�un5����~؄+-��
��r�j㉑N��E�ۘ�7q��bnT�;=^v˸:��Ȯ����b���l1ӣ#u9�����vJ�[9Pئ�sN�����u�퉰����x���w��Y%j�l�b�+o&[n_#
$�5�ݶ���dX䴴�y�	V��cm삆��B������ln�Ĥ�Y�p>�#/���c�����`RQݓ�쯵�,�,�c������$���O�I�Ep���I���5������/q	I�iuԼnln�~���j���,*����r�z�;��˯Z�F^�󺾊&���o�+oJ��V�&O�2_����p�ڿ�p՗ǇŬ�h��q_��Δ|�r�����X���ʡ4��-e5&��,����W������^E������uc'�偡&�/�����F�6����?m��d�^7��_�W����z�ػ��!�r����dQ���O;8��v�&Mr�v���ʅe��
?*���ӡJ�W\eĪM�^U	ٟ�g&�va��u��g��wq�ћ�;�ݻj^�>r�|��Aa�/�쾎�y�/�_.��tm_/������I־�5$e�z�4K��6��D�X��!�������U*��K#�߱������k6x]N槻e��r����/��Ҡ]����U2�m�D$�7���7����o�(j,�jd���[l�.ؾ�~?��d����M��"�v?��~S���x�	T7W~R�ߔ�7i��x�.IBU�e����ܥ	7d�c�m��D<����o��B�%Q��M����䅁ŋ�ȶ���$������S&���`��s�z���(n�W�Y*��`qekY/%bh���er����FH�䭜�!���l�B��b)���V����l�6r�W_��r�s���ET��}[���֦�ui��5������&��X��,��j���e���f9=��_[)y��}&�e��\�.z���BNO��"�j�"��+�'+���ы�7�+�P�J�ZU���d�J�+���8e��|���������E����S[v(&G�D%���*�S[���ubm��dm�ϴ$�	�_�gX���\�ķ�gXvAg�t��˴����++��v6����jY��ו��K%�~�L_>˿ۃc(p�g�J[�ֈ��g�����e�~/�E)B���k�5_�̄�K�TV2����R�������X\H��%�?%U������KZ,p��M�S�\(�ڵ"�"	pc0<�i����ݮ):&�����X������/��
��"�P �1J����S��8z�$�LZ;
���v�h���#Q�K�ˬ~M|�2�iv<�~sZ<�lif��0��섅jaT�m��*sXj�f�$S���5�����w{��rB�u�}휍��`�k;-����b�M@������s-Ł(dj�x�c���D�y�����#�?_'��?�R�ݦ�/��S��i��-�a�Ae�a%	V�Ƿ{@�{m����{�ɲ��U�5��7Z�m��/K4���ts����ZRy+V6?_�,�f���V2}��ܤ��aW������Tc���|�	�����'�������6l�6k��`�n�S�/V��֊KN�q����w�=o�¢K��-U�E.���nE��a����E���X�I�(����i=������+�~a9�@㗵}\w`�!5������dgX��=n"z���/��\)u�g/��;�X����]4	�q��>
�"���ςH��ӮRz�l��0S�/|&�t�2���{.��-���c�`s���a�g'䳫I�B����,�ܑFG��4�	 �"Z8�p"��?�����Uʷ��ip��B�q��KѳϧB�{u�{u�U���xE�؝��\\~��۱��6��˕�/+�;�ɣh�\%�㢗��ޫv�v����I����)|:�aN�uTe�pή:7sU�cq_�6&��^u~��������"���<�Yd��ѻ��@��B����K����
��a٣���!n�[�Zo+���҅gc%Q�=�\��+�۝���Y�JY�:hl�����ݎ�Y*���B����CM�Ò��m��>��$_Se�d�l�6˽��]��/����R�-��%���r/ʶ�rv]ejە��Y},L{e��oi�=��k���r4;e��lk0	S$JKt����^��F���Sn��)Z��:��5�c;]��ju,]F�[�1rV�^H��6�|^�W;Y��jueF����]�k��;cc��eQ��+Iګ}[��y㉁��g�ubz�U���>k�#s�%����O���ť�&\N��]Y
g(D �{z-���DM��������³���&�'��ʥۻ�2}d~R�ҡT?j!'�ۏ�u���2�,oơR{�+W�)Fe��r\����φ6=�筏���p<�X8��I+��M��?%�Y���f���&�H�<�v4�R�P
�:K�mYnV���e-����2�]���D��Ձ�bU/�J�0j�n�<�$�����.�o�Y�kU}��=�v�^�'XQ�#��g��`i۞e/˻�ir\�726��OV���Kv{���{"V�R�䕓�dCt�M�����ĳ��w�ڣ&돲��ܚ^O��hK�k���fb�_�����M��h�K$Z��ߚ�n��_����-�dh��Fݪ|C���Ce�.u��'�Y�߱�eW�sf1���%ʥ��՟;�.h�U�^���e�ȠH�Ģcga&��F��rn�l+�g�r�� b��}6��ŖM���\V#gɢ2R�������+lf���g ���4Ci+��.�@��J������q�njҥg���B�����=g�+�'�gȱ��VN��݈`�7��l*�6���O���RP,k�̉CKw�� ʫ�`~ơ:����)g���l��n�R_�;8F�,j�}F}g�@��}���Z�A,�U�eR{PQ�����X���it����f���O�^]�ntR�j��k��K�2�d������椕Xɴ�WtQ����_��u��|�޾�u��ss��	�J�X�@�@��K��Ï�k�(ߚ���UN�[�ѫ;��̣��9_����F.&"I��V5dR�x�{�v����4��yx+M8��ig>�N"P�K¥��%��	V��rϋ�u��FQ\i?�������_Ieկ�rI�;�,�$�ۻ�M�Su2Uo-���ӣdRnq�2}�)�X�ga[<�n�R���Z����j�SwY(ik2Z��BEH�EV7Ϝ�ĺ�t�:7��9|4q浣�l�tK�㫚uIr�Ev��uWo�EV�:��qj2
�W���N��I�6Y�~�$[�l�f����JR�%��>�	M���vm6lGw7�/%-��P�-n��^�EGe�̇������|���H�]m?�]�q�=�����
/��o$�w���(8�vH����˞+�㫙_�tS����~���7��ټ����ټ��7/A�?{���S6�z����mN���~N��E}��vC��\�;e$q��9��o!���7c� ���\�;M#Yu��Kg-�d�:T���+#Yi��l�l��|�HY�6R��r��t?ʕKn�]���[��ΖK/ɕ䔲��&M
�ճ�F�U�R\iR./Qc�F�������|L�[�������8�(�T����_�x�8h���K8�̋N�5�DddCK?;m���
L1�]���B����r��E�&��[q�3�u1�ȯ����D�7�l�����nG8�����a��Ukˌz͸L^��ԫ�l+"
��曹������ɥ*l�D~�'������[����0a5�nUʟ��@�y9�v�wV0Y2��e�S�/ ��gZn?�Yi�/�_M�BYnO��Vl�&��B�Rac>ᤧq0<��w"a�O8o�:7Y��?�`hR,3�}�����_��^6P�sUς��¡�U՝��	w���'�iJ�.K	sD*DՂI�#(�6�&�����r(.|X�:Vl:�Ⱦ��	=YC����'8������]��ϻ(K*�V-���ոHu��P �6��Z�ςFZg�;,V�Uq��_?8?����,���Iw��m�&)\��,,`�65d�������+���퉬K#e���i��݅k�ZY�35���Ly)f
��a�"��i"�q@���ֿXnE���a��S��^�nӆY��IY��<6Yɗ��j<��l_���$t�r�µ�\��ԡ*�k�ϗǯ�~�c���o�]�K��{<������I�>�I���#~�V7ȣVK�|JY��H��q3����"�cIv2OWn�"�dFI��J�#a<�(��V�c����~5��q���p�����Z7�UZN���M��Fi����K�n�'"ד]�EuWD���+�Б��k�9��;��P��d�jH*HO���$ԐU�Uy�a%�ˤ��Tjݗ�V�:7㽘�v�~<�>n;#8v��;��mԟB�
&]h̖rI�;+��g�
B���HTb&�m%7^U!m��u��ؿޤ�B_�ǭ~��̈́���Ȃ��_	 ���$�f#�ܚ��勶±t��'g6�����J�l-����w%���kt͊O��nFv�#k�)�����Y�:�s�I��,�׻	Վ��a^]��՗Q�Q�����W5�J%҉E|�xo���Ug���~���?<�ל����6�E��_�e���'�b��5�d_Q!좜jl��bd:ݿ�A��}�j�!S>,"��M���މK���ߵ�ըw�����&���CD�|�9e��l��|7%L�z#����l�~�ǋk�xk�.>P���j�)��ό�]���^4������K[�Ҷ[�W2E�S!�+k+mԾ_QA���܎�Ws�)�kiY��;��b��ƃdk����fZ�Ɔ�+Q|��r��nT�D7$\�y=)aɲ�ir���	n���j_�>���(L����Bi�5�m��[a�nBҭ�b�l�n�_>���E�J�����0��'U��:���.�wj��QQ�/�6	/w��h�N��Vy�f�*�r�o�S�a4���ܤ�r��@iF,�߯�K9�ܱDߚ�ٿ!�w�8��rH:�{��������//�I��l��:�jY��`y�"�k��q�,��`�vXsҌ�"���>)dl���!V"wu����5�l�7�{{(�ذ���Z�5w%I��k#�_�v&Fʷ!,h۩e�-LBE-�����E���Rm�qk8������������	����$lC2�'7[��Vp��%���ӫ�]�q���I��]z���gɥ�aiE���fE;w�R߯���ۤXQH��֑�I*��ȓhBH*+�������Y7�=o�`D��G��V��z�a7%�Z��=�i,+���[��[�lk��l:,p�nI�^q{�q|+����eW��,񽔏�b	�mϒ�t�V�ݽ��de��|��]y�)7!.RV���g��_�����xe��-Ye�6{��z��I�U|��n�o��Wd"&�����_"�x���*�L��b��mb�����@��oȗ��n�m;dR�|�˃@���F�b7$�*���6'#ie�������k8���4c�
v��V{Q�7l�Y�c'�ɭH���i.�XѕY�W���\}y�Qhh���bl���%ł��"U�%e܆�Y��ǡagq,ұ��B9��[��^�5y���5��c?ߎ^�l8z������:��ڂ�;���|�ڲ���-Q�F�wḵ������%V,ix,k��g/�����dVl����k�!#?���hƼ���ʥ��M�7��i��M"�q?��xpa3FڣW��өvƝ�Ų�I�+�m�q�w^���c/�U�E�O~G�yK�k�j�u�qg�X䍅g�ܯ�
���J^�I&�F\vV��*A��5�66X��\Y�k+���2U�Wi!e?QMy

�Yd/F��iWv��=�j�d&���Umy�M<2�Whѵ�_6�5q�:���ٮ�L��U%����E]/����U��/�덟����u�kW(l�[�,T�@��vqI%S��R�w�[n���JYkW<�wݲ��~��Hu�K���N����7*���ⰼW��m�f�ke��%Y��G��θ�T�������g·��uܗ�|A�}/���lW�\���W�\۩}k�PqX_y��b��NwK����m*GR��}*)��w?�z���~?r��$|A����C��NS{���*��Ei��W/K����QR�{ht��$E+\�{��X�\JR&�;!H;u���M����I�>��XH��_�,%�7��/��Y{�SK���W�������玮kWmKߎ_7�}i!-Bs����dm��*�זo��eiіݴ�5��;��G&��Y��O,��7�m#���ɫ\���v&���Ԣ�o�J������V"�r����03��$�ʒ����f�}J�#(�
n޾J!�ewd���.��)V>Ȭj��/�3"M�@�F�W�m�l�}�l���5�x�2E�&J�`��p��?��H�*L2������7%z
�7ZƼ��an�I��X�AX�F��*_*���K�V�7a6��Q6��I�Y��4K9��¤�Ԋ�&O
��IW5$��T"�2��m�ѫ���Q��K�\%���9�]�bY�6D#�IE�H�sY�j�����54�)c	|d��,�J��iK�q�x���f�a|*2�!b�Z��݁J���;5���:}$��>���*�K��T%;ge�_�����h��_��W�q,��-x--x,��,�N)^EM�ǿ��?	M���׷j����"L��_�׿{�/�$W�!������\���ݔ�ň�XB���Z���"�*�J��;on�����.��L�����,?#jר-��ܫW��'KE�wZXV�O�^κ�`�Z ������7���|?�-�d��O_/��FD��|;��0���B��~P,�(|�l�HD�d�^���_�>?�jʼ����q�8����,)J��b��8p�f��T�vtqớ
������o�6b�w��f5����
�jw�mFh����7)W�O�yգ���<<�.-uƽ���֓]�}�f�7_��\�<�ꪸ���D5\�l��2+n�[?/�Q2�
69�HE���&ۥ�/�a[�V������6]c��r�2��?_h����W=+g8��V�';��;X��JY�-����͎K�l��0~�V�c�������5���|R+n'cۖ��R_�#E6�"�~%����	W�V<+R�WoK�U�_uv�\y�s���5\6���vk��.�J���o���;Wo�/8o8���̓`��K!�ޯݗ+V�]�KR߶��-�l��?M��$jJF��J^�͍?S����)S!�J�1����-Ծ��R�i��;Q��^4����:��WlW���3�O�q���w9�W���÷�Z����^��>��/��~�x�@��� ����+����8���V~2v�WS�V��ܕL�k-���.�S�+�J�-�!d��e�P��1$�|yF)+<1�Y��Exd?�����	Y��B�$���c��[���"���Kt�5y@�%�5�k�*�U��W��G�|>��n������ψK���V�k�L8�hݵ/�5�xo(��^�k�4h�	������͆�kTq�Y�ѫ�?�e�濜�|N���Q�����p�������kJ������������_+-��-,��Q<|�n�֟S�k�9+���v��BOaʠaᰂ�g¤�M&W������oK46Ywv�l���J�o�E%���Ϋ�)T�KoWg[��+���4���*R�������%�D%\�=���w2�<���K�&D]X�~�$��2�݌~♈��k<�d�ʒ�K��"��ak	.fU�͆M��I���V�Aw?{M�e�r[��F�-��@���3H��ݗ���Y�v�"ƮiT9fo:_V5RkQ�.J���i{>��6�l�y��J�-�&��}�	`\\H[�z֛v牕[���<\m3%�!���%|��"�J�5`g&��]��IM�ѻj���l+!"�@���Z�uc40����r�8c7��wi?����\n��Ȼ)���C+��
�K5��Q:�]|KKD*E�
�M*��p�c~�V[�ϴ�����P.$hU������>E%p�e�y.<��	�"��cW�_�n63n3ο�M��0�,��C{��v��,q����^�gG>H+?�H-���]n �+vy�.(͸ˌѺ�l� �$Y�`��Rx����ȱ�,�I��T�r%��Vz96�x�k���T^E|�hE�7;Z�گ�ߥ��K^&	����%�y����V�GY?��mO��5����ӗ����z��tK��V|�h.���-�8�l`�Xa3�AD�X�v���v@���	�2M	cW���Wڻ�7�����Mv^�֓&^���ʷ2:����Y�µX�5��R/(K�K��ݍ͚U�^����_������{��e'T��W��@�ґI�7h� s�L�?�[�gd��4+^'�X�\*�I�9T��#e����<���������<6�X��f���z/�j��5����6�����с'�)ܔ�o�V1=dU��R)<��^��B��y�K�_5�j�͎��fяF�ޝ��](�Wp�}��y��ۆ�(=w0ba�+�R~}�Z"���D7�ǻݫ���̌�__i��z+Zڝ/' ����/�l�whx�7�]��q�����+V������s�?r�{��x�Ta�.�G���^��9z>Ht9Y�(bKE �bC���n�+(0:�C�+1���T��-�x��L��V�s��P��k���M*�B�q��"@��x��[-���ke������-�v4��»���jr�;nv�e�R�-������98w�ݵ��jw)g���1(���3s�q6���Ც�[+Y��[u/8<��v�V3_�����y�jн:�e�h����dOX�I{��mK�ǆ�5Wf���Ū=m]�â7�~�d������g���HQ{8��&��ǊT�/��YFO��SM�ݰ������ݦ�2!���"�C���rJ�V"�����*����,�rX��;n��[��km��xl,l��6kh��Fi݄��E�ggH���JY�!B����C���{�|[�_ZƼ�J� ��H�ќVp��D�Բ
O�h"m:�o͑�y��&�[�H�����;�̷ߕ�e�v���w���1�F��a�.D�Á�	F�;Q��Rf@�zK���0:�L&e[x�t.FA}-�uF��ʑ"ћ"�|c1��Sm�Mܗ�ʣ%.��FK�ȂùaI��n���QM��O�ʈ7�[���W/�V�e���d��,��K�6�;[u��T���y�'%�lFc��ڲ-�<���E�_?�"��X�I�_��)�N���I����v����'�s�5�Ţ�~�iٟ#P0�Rm{�-/�H�?�g����)X��x`���y����I)\���݉��'�I\:�hl�˹�v3X-�����J6!I���������K���qu\*5�NO�5���g[�F�r+�-~|1�p-U�U��K���2%,��p�}Y�, R�	{��O0�K<q��0q�Ԋ�g���sK/�I�w�~�<�F�Ղ��	z��7D��8,�a0��5�tQ].��v_8j�L���Rh�����4�㰸���w������Iڻ��m��v���#:ၵIgc�۹_�,���tq��K��:14��c �����p�<2�ݽ/j�����'�"���ݯ��b�\/�̂��M�U�V'o"ּ���Yb]T�E�����c>�c^����8�pW)����J!�%E�zNL���~�*o%~/��Q�����k:ε��w){��Hyz��*����cW[%s��ܵ.N��{���Sr+�]7�A���ʥ������?
E'��2���n������£u}۸mK��F�:�maǍvk���E:��o�j������'6k�����FS%��x{�l|���*���mCaTiնCJ壒
�����&ܰ�[r#���T��M�@�a�	g�r��a�!I�2V{�T�vJ��E�0)ې��巻�Œ���s����k�e_:U|�f���	�G��VO��M������r'��\�Ֆ_v7F��0�����c1�WW�on����'�nI�7��2,���(VVOr��d[cr-��.Ko+r?��߲�n�I&K�]���lfl(H֊H-Z��R��<V�e_򨄃����w?-��,}�n�F���/����[��i>�F��r�nڗ�j]vj+����j�<ў~Ȭq�u�����~vb$����4�'��
]U��m9%
&]"�Ռ��_�?؅H���l�C�߽�j%�̕'��j�%�nQ���.�!&�mҵe쁒�X鲦��\2~��y,�U��4_q�N���V�JM�6����,�e(lܛD]���=&/}�,����њM���
ܕE����-*om�?Y|���X�������杸��F!��;
J[�~T���Zz�o����1.��´�V���	4��~�&���M�h�z�ir��2\�M�,�`�nF��D�&=���e�$e�maj��dP1<�/�rj:�mL~[��z,�e-�^��4_z�g��_@�,�a��W"a.�6�3��$l��˷e����p��D��Y����q��c�E�ۃ&���>V�~H%�^�	d6M�'��ɛ|��Ѷ�(�GB����U��6����_rw.��z��>����ጣ�����Ν�I%ru�ʠc�2,�$�A�����Y
�h�h�ۂ��}�䉻g.�U܁�����۔%bD�̰\k���Ȱk0��1�}O%&�o���/������B@��Z%V�PP)��~���~i>=]�f��!H����丳�e�D7;e�����k噳h�â�ۉ��MZO�)<J^wp�kZ1��U2e���zˮ/\^�K�\@�AU��?6��sa�U�
�Z*���Y|�7�{9Vޗ�dl���yᝫ�㢢�����H��c]�����k�v��/O���'�۔�qȮ�e���%�5be��Z�o4e�Q�V?V?P9���Ddh���Tn���f��~|�WVE���*ն�caY�fj9���ܯզ�kӹ6�zƣ;���D#��,E�g�����k6�y�͕v�G>6����%X�ۺՑ\p�K�`Iῑ���dR|�Kl^
O^�Y�*�	>xٰ�*߆�z*�̗�����ї�;�S�wn��D�Q_uF����/��\tXos�BfX��ɟ  kr���"���J��U؇�!c���~�p�N���V܋��[�e�)�hN��d����H���_i!�w�XV�����u��wv������n��ŋ�qYv���ZÊPې��Ǌ����6�{N*�+���ߦ�xd��/�ۏ�!�]�^B��S����%jdl��KR�|��,�W����˃5��>~�+��Hըv[gLҹSleQMN��Gi{,�/-���NVe�?vҳ�e�r}�7v/I*\}��5����a�;:G�=�+������.Wg���u�m�p)ΎluscM<2�h���6�2^�2���գ�
�Լ��F�;P���y�aV7���M[�n�rX2������L��O�\gU�'���e&��G^L����\�c!�'��Yl5�<L�腐�V���&�ߓ�۱��Y�ۥV��	����*I�7#,)�)=onMN�ܓhȰRu�֓��v��_��q�c,�v4	&�r�b7=�U��7)5%;n�?�q�KX�L�Yc��T�@��jʣ.ʩ/Ҥ�Ҥ��q�ɩ)�[{I�dk_�>���?g�(�n��o������ck����?�E��rrU+���[Q�Z�0�Iv8J�z�N�4�_�e^Vw˨˨�LkD�W�f#j�ۖ1�8Ѹn5�1�R%�9�2$�*ĽcU�`��ݤ���ȄXZ�gqk�	��I�"�,��Z0��^Q�=V7������"p���E��^'���c7�Ul'���˵���&�B�u=o&&B��%6E��c'��ʤ�o]�J�59�oֲM���Z�@���|y��aPL�.O��g��X���}��sP$W-�7� ��Rұ퐸u�	=EN�Sc��mo�M���h��[���p�j+y�(��n>��5orRݳ�I��ZX���I����5$B�^��
�g¨p�>��gf�ۖ��~Bݬb7�����87mXK�D���������j����۱��I'�a���f�s�QZ����Z+�{�u���gV^��7�
7���q&�q��&��H���Փ\XB.�P�0�0Z3@��ʩ9�\f�����3��N}i!:��]_��^}~���K.!<���5s@�&ͣ�3K����K���~MvY�r������Z���!p�����#P\�s>�u�/�G��㗫��^�ؘ+T��dR.(�bÊ��nM"��rV�F�*�_�⒨���n�R���y���d�Xc��+��(��~/����۳�"��Cv��Áe��D8c8nH���05���P��~�a�j�@�F��c�Z��<�z�D�߆��˯��Fwh�&oQ(�Wh�՜��mQ���������M�������ϋ^Ua���_�����2Ym��d�Q:\��7vJ�V�!R��~B�j*~ڌ��k)Y�e/L��=�Ƕ)Ŧ�����*������}�v�ݠ�7<�%e⚚ƶ+b`;'�6����24M��S��F�'����J��yߕO-��u���vC�d-l�E�w���������Z�ȖvV08����moc[���+)��X�HqM����G�V�Ʋ��[�Y"���ev<_vߟ�h����X�ԗU�h�I�<v��R�zn�nvB�S���.Jo*����Yq�����sa^]�/V��=a4B@�ͅV���߆��jߎ���j�Ç��08����@�J��_��_V�_q�"�וyՕK�)��B�Rm܄���w�8p ����}.�[r5���f�M\K{/u*ۓ�\o������,qR@�[�oˌ���v�R�[)��f�W%ßIײEIë�*�&����ն����ɨ�%Q�5�X����v����*Ҍ���]ݯ��&���7,E74���qv傑A>�K!4\�n�׫���%_y�Ȗ4YQ�BO������YNյ����|��J�lD6�;K.%R�AUur��Ȝ*�,�«z��;︻[���c41���~4����nʼ�e��?�Ղ�a<�}���O$���w�.3qW�]U��PM�M��*��������g�vR>̣͌��gVE���7R�Q��n�)	<���g ��Ȥ����kJ�Rb�1���m��`��������-��n�`la�(�:��&���E�ܦ����MM�>�#fۻ9J7�D���005�18�,u��ܵ�M��}���V0%����01�.턅�cX�I��v]|��1?�<�����vU��%���r�+�:���*���)�PZ���f���
�*��v`�t�;��-���F�BM��I���U��w��)qE󿚲�]�J2z4|��dY����"ã>����*�a�߱��@���w��8y�y����[���<��Xh�̺]N�5��g}٦Ns���z�gX��7��=�nDM���a9���@㵢�|k?����s�=tD����5���B@���D$�U]U�&�2�j���.�� �]�sF]K1��x�+�wbi$��+7e��&��}�N��O�T�~�D�ȳ�'�:��˗f|^!�e���d�f����jr����P7q��=yK�!����dBS�/�_�&�
�.V^ܭ�V���?r��ncȯ���'�n���Z���ܷt�
��ڱ�WJ�tRF3a��5�-/%�����I�F��9��_5�Ѣ���o�Fto�R�E:��o�j�\te�U]-_|&�M�YGVY~}=|X.x��bU��ϳ���.U�BA�����H8=��9<l����d>6�'R�d�^�t�����*}ceQ䔫_�io��wm��ʙV�1X�J;�N����#eRw"A��gdnM3�;������슁����X�nܡ�׶�eQN�_e�@�`�i����c�����iK72�ݕ�%�i�7;n��M��bZ|od��۲���b8nV��T�/o�cc խ�2-�8n�����d�E/Y$~��J_eoѢO����jT���O���-XU��;���r����P�²Yy%�V/���ڍ�Nk�sז������R�9z3���;���藿�ї����ļZ�񙴬��H�h��7T�o��RA ��Wc>щ��l3c��j^N�V;3��!n6�5c����Fn�F�V��+o�e�����������^귞��Y�����,�ݳѥ'��n�v+/��/_�W̪�D���u�g"���a[ۓ�b�����cV�_kvE'�p������'"�Fhu��.��.*�:�0���^~�+vg�/����h�ٷ~�	V6�2��������\H�3Y�X�AQX�a%�Nq�,z��c%��Ȅ��XB�V��J�l���5��Ԝ�T�ac�}�[wT����(�d�:5�?�`�ܰRaAQH���#q�.3I���].a?��^�;��f�;�h�%Z"aQ����$��h���rdk��P��lw)g�+�3e@�X�7tfϣ*�뫡́I����sw�^�\�?���ҵr�m�m�W�%@�u�iY*MgL�큂���ϣ,���m7%��5k�2���́V7+�I����2�[f_?e����vإ�Rʷ��%�n7!/�Qǿ����j�*����,-rD��_Rm��_ʛa[�����	���YV�"���
OF�r
���U�,�VEkd�T����KX�'�G��^�\�W12�q�����zї��w5�|�n:�/}٨�:�o���ޫF�u����`D�� tdFK��K��W��Xr�����Wﺗ�}�Y��	��M��S�K�b|脁Kݗ��W�5�[碪�&Γn�âO�^��Ç��ld+�%�x/�NV�#gq¤X�R(J޿�nzU��?蒫�,�v�
O	I*���W�\n�`Өf"/��H��	e���ݔ'�}��K4ݲwe��H�����)Bv�o�qv�e/r�f�J���	Vޣ�J���u�w�:���"�8��f�������"��"����Ob�����߫��xk��a$��0�1��y��V���ѣ//v�Z2�p��:7ΩD�UO�ڻww��w5V;���TW�YU����|�v�Ӭ�<0�͞��~ܼ�VO�X�#��G����M�[��.�ij'�3����ʙ�풣�^�!����t;.¥������+n��*t�L��)���jO�����nRW�[-w�%Y�m%�o*��m��n��R��S�m����w*o����k��1z�}�/�����L_�)M�����6�"ݝ�!�5g�c���o���o�$H[J;iA�Ex�*VnYr�(������r�>���d��|FOk�N�@��d��Y>�o�&�8�R�6���m�K7m�2�^?�Z�W��P��&�_����Iyu��x�^�6>p��㴙F���U���5e�Ỏ�^wsU��ۋRx�?��b!r��T�7'�w�RZ��!<�IaŹg,�,�������dѕeQ�����ukD�r� �j���<�.ǻ[`fqF@��z�W+d4_=*��ʋ�l��J�%�Q6�`F��ȵ*�������}בAjɳK ��;�+���nK8�Rn����.�H��H��T��l'�x.L�؆�+����0�z�~��c��&��ݐ�6���g�w앸݁�!d5n8h��U4R�GY�o���h�mn5c�O�&�34&�)nk�eS���J9�$.$�C~�5cV��%��U/��1�jE����69=�A���b{pn9$��kZ�бЂ��EI�'�Yc�&��́_'��IX2��^���s%�+�g�#5���Ŭ�J�jFDC_WJMف�&�r�u��ܨ}���J�u�}��X�u�����갺�c��I�ɰ�H��[dY,����݂���d,
�Oe�?,D��.%��02����Mm�V�M���m���nS��T6H�����2\V2����B5n�2��0��;��{���X��r�߂��,B�tS��� ��&�f�'/��y�?�ѫ�*�RXK����`�K4���~�I�Wi/����	�Ϗ�b8��&�e�K�J��n�%��G�%�K�Xj�(�u�q���ƿD֊�:*���q�ժ7o/'5Z7᪵z�T�V���:����u�<�h�|�z_Z��p��Ej&�?���	t�0�j4}'��&*���ij�����ϓV�'��
Mհ�d%���h�D�B�R�+��Jߵ�nR7`��69�T�S@�mϓ��,v�R��k���&G>,|�;iJ����ɢ��,\^?S����v{�ߛ.�?�>���X��s�P����/���B}�����]aX?��-��Oذ��#w����Nx�~ڍ�*�o��٪���,7�p���EXk��Ͼc`�h��Q�wn����ѻV�8mZ�v��h�T��^l7���}�to�u/5R^s�V���~��ޗ���&�� �h��z��d�N��������]���+�J�[��������+�_����D>�H4����iR?J�V�{,����~J�R��S5���N�)_�!\R~K5����*A��rYM.N&�v���J_����ʁ(d�+d����I��ڞqQ�q�	'gé�i��]mF۲��^�f����V���U1�^�������-�VC�B��AW~B��c�Ʀ���Px
���Ts�}���S)x�����C��DA�Hռ�~������S�ը�q��[=���?���2�}�n�gL�g«k�W޼��	V�eZ7q�U�~���M:7��WG�j,~tvo�R`����Z���g'��H��}D��c�����ȕ(�a�a����jIe|�JD�zUc)D!(P<6x9ؾ��P��)�l���fw�W��&qX@�\�oD��P�J�9�����t��w04J�tJ��3�7)T����o?�E��H�+<�&�zǬ���ò��7����Q�}�Cn_w04J�^e�Wɿɩܖ0�/�y��`l~ܡ�9��HJ9��)5gvB�vK(�4.^k钅�#+'��}���k
�i��p����|�F]�Ejmg	��n������0<��%P7�s��v�qIВ�u���:�(��[�+b
^�����o���-+�pHۄne�8+��4��]�>�vP�cݯY�����,��j+P�h�W��]aIc�&��]�%P4J\��\�-�-�~ғ�վOX�qenQ�����a�F�'8&���I��B�0)*�QdK��pk�(�v�����EF�W�����]}�,��շ�U��B�x�*�5/r���K1��._]�+���8)K_4B����k$M���R���U�I��aT��F>�)=�2z/�r)z�/�}�M�����
����vAiqX��RF`\c�}���17���g��7l>ʿт��IvU�͟\Ԓ�|������2Y��o<p4`~���4���֋t�Mv��ڣv^��5n���ݺ�t���nvp_��!5���u���Z�9z*+�ˮ�f�дK��u�_�uuj���E�����'�Y����	�/w4g���T�s?5|%����+�r#{pe���T�ۏn�&ǎ"�!ns����w�Xk�5�WZv�K�Y���a'�������k��ձ��qIVXN-.N#�/���b%��K?/%s������j�,mXV.RjwCg�ܒ�|��\_Ѧ���AV�����OMa%D%X��gn}<&D����m�dV(���u�n2$L�TK�+�j7�a�^x�,c c>��ޣz���;�o�F^^_�z�o�Ev�/4��f�z��y��:�5g/��<���1��לlM��c{7i76�7y4���˕�����S�ņ����YvR52�#��̦��K��{͌���[�����$wv����=�l�*�%��_�����kW8V�)� �d�e�%H�Vv����i��E�A��dn�C��Ɉ��X�l���edl_*ݝ�Tv�6[�A�m%�.W)!e�\��{a-�:�+��|Sv���*����)����F���=xV�����[��ܖ�Y�/�����+?��ʭo66��*���ۿV]�w�P��vREcYY䐶pܯʷ���7!����N��S�8��k~A��~I_p?%���J�x�6|%���R�2i~z1��U��~֪ڗL�9��\k�sU�g����z����dݚ\�)0��c�I�7%�i��n���,q���2�>e���ˠ��m�Q���jE�I��!�.Q�W<F��Y/ ���P��ܟ�6厷��%���
��*�y�jY�M}���x)�\yϓ�S�+���dЭM����>��_5I�	j������%�^p��BUI�y��?�`ݰ���u�ϖRp��R+�4���#Y_ݭ��6Y	��ӳ��^GKi!��^O�_?��~ګ���ߚ��J�h�k��w$ϸQ8h��/Z�.�I���MۥV�ᘁf�dB7c1ӵ�1|0_�6q04�o�ZZ��&�j�!ZW)J����%(j\�uBp���ș��j�c�Sb{Y�8��,9�Q:�۔+%ݐ�/��`y�gc����E,ϰ���g/��I��D�;d&�s�����?��!��ɹ����=�|S:�Ry�RiJ��(H���oVn��d������l_��(j�ጸ�W�K�I�!���-�o���8n�ڲ�b�yz��>�c�#�����
�*���!%^r����_�ߌ��������a����c�I��t�/���.�!I�u���4���?�� ��Yګ�ρ���&���^�U	c���~g��;�*��7���_&b\�\W�ՉՅdD��U��z��������k���ma�v�;�}�/UD�ͣ=n1�ц_Z7ݘ��wtXB@����u�'��^�c�;US.��a�ϯ��2��k�Ό��k��%�?�e�-c��
&E��"�����<�a$Ԗ|ZV�-=W����ݰW�BO�7J2��v�'��n߿`܉du��'���Q��F�����"�JI���w2�V��!Y�,�Iz���Rݬ�`�\?d-��C��|$7W�c%X��eT�i���Y`�3���iA%���,�!Y���ަA���;vRV��r�ك�JE���&s�=|��_�^�r�wX����
^j�Wf�5����۴hѫ/F����]�U0͆l3Z�D��E�^���Z���<�����ׯ���|�5�}�g���s��Lm_�`�R�>���Ur����C%����&�o�g��5��z�F䃁�M�Ϗ�J��V\�l�v�r�b7�n-�B巋�׭�q=Nʟ��,�Qx�H�J�6���Svy�������cr�Ȇ�ʨ������ՅguaY����^⿆?��|��-(VUj�싇^%rV5�|^�^�I�с	g�����_��Ѫ��Z�h����a�8��9����Lk1�R}�ƔC%��!I�i����%�%&|�?��$e�9y�y2����`��V�j������F��]뤼��/�F�
U��6�Uf�̌����RFU����⯹mᱤ�c,�ߤ��QK�u@ˢp�ݓ�D5ബe���ۖvbq:Ⱦis���	%B�°h�X�Cui%U$�
���ѥ'�,��'��:�_�O�^�	���{x����Ȳ�\rd,z� q���:'a�3�����$�74��2�񖸤��R�]����V�k���kR��5xl�����!,�M�r�e+~z�[Ϋ捗��*̓�1���a(�Y�`pm���~�!�����r+�"`W��t�9�+D��d���2Y���¿1�лa�/��E�����Bm�b-�,B�\��7�4d�lCv���,���V���,^�J���X�g�P5sG�9�wn�������By�H�.0w#)2!08��-Y>k�?�p�As��Rҍ��"�,�[�\[_�=o&m����q��Wܵ��,�'�2�J�m����(U|��������c�۸��h��Y���O+�Y���i@�?�w1��\��=6�%nT�B�����$^�6˟��j�+X����;�cp�F$X]H'>�N��nPS܄dh��ɵ�0�	Cr����$O��'��K$���������rR`���Q������e��߇���8�'|�h�c3/�a������+�I�?4z�.ZQ�:8ӗUƫ�¿D�i:�����������Fiz7S&Ns�v�5g���tRy�aF�e�n�=q��ƙEI	"ґK3��,�j���6���1��P7sU^L�v�<=~�����߶��m\�)5&h��19����v�f<2h���sAUAQ����\��u~�|�����}��͟_,��(ް���~vJ�֤lfw̃N�([d�I+sʌ�;tP09�p[��w�5��&���\�)
A�~oѓ�aϤI�@�%XX���i+/EJ���H{��4�B��V? a\]y5��v_�j��R�ʤ�"`V�U0�;Wg/EV���f��Ns���Ѿ��uv�T�0͆l3](��c��5[�ўk�{��ty�U���Dm��\(��͚ϳ���͚0�\n���Ԃ����{������:�df�־E��ǈ�uQ���Eg�"�h���U�@��u���������7l��Ш�T~�V��Y�	"�J��z�#�%,ܦ�Y�X��t�e.�e �x�VSc���$h��aA��~��{��Tdv��++�7[����G#T�U���
��#E2^ڜ�ʦ`���]�;S����2;e/�c���²��|�.��hݫ��;�(������ޙvi��v^����|�����K&���k�3����K$Ո����<&F�V<�����VR����_�BaJ���g2�2��^�����ژ�$����Ϯ䞒!����}��Q���&��I�Ev�˝t���8�Z�4ؾ�R��4u��?�;�+����M7�3��Uzܤ�Q*��00��*��U��rL�泂AURZ��G�h�&����"�~!R�o#�?q�����3,mK)������J��޺]O�d�b�֪ZHE����q}�2ә��f1��yߚ
әh����͑���uc����,�k�-Z�u���e�
���G'D�r��q&�,�k�P5����(�|+w��eR��-�-I�唚�9�0�`�}�V�7����&|&n�:���ԅ$YW(ܼ�4Q��IN҉�y��"߯����Y.�Nί�l��J�������SY|\��¾6H���
U�J��!g��s��T�o�-��HR)��[�7(J�+r�;r�N�Q�F�܄͹W�􌿞������<��<��#!�10�'��l���%�����Vv�J�}݂�܉�׉���#�;Tݵ	W��q���(����Q�Z��۸���	~?��`of0���Z�/����(�%���q�6��7�7\v�իv���ݝ\8e�f^���:%��Ḥ���M��^y�n9��.�U&��a�_��%˩ڻGD��tmuǎ5�e�ᾭ�ӣ}5SFI��\]�W-�:��e%~��Y��	gv&���5���j�A_g���D����/��?v��{+��_��D�p�V3׳���>��~��v�ov{�=��l+Cos�����Q��E��Fb�qµ`����T�@����ؽ�7�?%mù_�ʦܹR
M�_��;�w~*=�}��B����o�B�0k޲)<���I�M�g�6����oQ(���ѽvs��2i�wݝ�}҉T�%�3a��Ev������2����g��d�U��d�$�M&�I�x�����;ܖ�'&ܬdp�V]7�!N�q~b�kiC-��l��Q|��g$f+n�'��Xn��\�r;l5bm����JP�S8k{*M(�ʱ���^��n�/��~Jەo�X�bu��R����a��T��)|��)�!��Z�6�Kn����b����Y��mӶq	Ca��[�{}oS#Yv���w'�e����\���J�%j!���qݶB��S��yJ�\S}zwv穎�̜?���x�B����5-�����{�c�K���
�}�B����ʢ}����[�r���N���$�O���}�\s����ɨջF���6���Fxo��<*%&��[�Fo��S��l�$6�M"��ϵa_}��m�Z��Y�]�Y�{����X֗�����D�A_V���ݐ�����r��*��iX~g�pʴvI�jUc�&��&�gI�Oq�'�,�����בU���"��!B�YXm��y;"���XV�k��I�j�*�������[��W��n{?����܊�BT�`���+{��2)E�Nτ�/���o�\S�����i4J�p��D����VuK�>n"a:�����y�K�/.��5e�U�j�
����.<�F!*��L&d�_1�c$Q4��`��*��FZX捋�X�w(ʠ��Xϵs`}D�aa���}YTg^R�E��vB��_ל�̽���/8w+��5lk|��K��LM[��̟6;P�����ƌ�yՕRiI�$В�p��l��FJ�Ϯ�a2�L�,W65r PKRm�Q��4�q��Ov�B��[�7� ���m���oW���Y��Ve	f�!�B���\Cd�V܊��M�⌶����,:�#%�3털�����}۰���m�.Փf�g�'�q�c��7F�O�*H��5�Cn��ľ��Xz]mYګ'��"ǆ��^2�UG��`h����}���Z7�*�a���G�y�n`nݸ��iW��2�yݵ��'<�0����U*�S�F��vs��2dӣz�uF��%��0�tQM�5�y���<7��E���Ľ�TIy�/Z�D��j^��S]�����=S}���nn��iJ�uuv�"e��+�.�'F&ל�܋n��"�'�v?�f\F�����g�u�/���,�/��|$7��+ ʴ҆F�%���c�Cd[e�wMcM��V�;�m��{�<]�J�זie���ܷ&K;'߈y�ύ�℅n�>7��{:�w���Z++����¶��++�R7��_�l�Yq	��k�*��V^�����E/4��vto���&M9�w�z���T�*�J+�����vwmh�q	�킯9~�?k�R�����^���n�aZ��ב\��o�m�l-�m��M��e��Ƶ)l���+a����[�^ƟN�H�Tݗe7Y� �Q|���BȠe%/��;e�X�H;J�7��rb�r+%�k2���Y���彭*�jrt?�+Q�%H҇��Ò�ȷ����_g"�JZ�L����b���F�H�R�����|�nKv/��u6�V��Hq�m����d��?O���W)Vd|���m$>�R�ֽ������ƻ�I�����H�-EO�]��;##�J�ҏ�p���*n#/m��z#$�w64y�Kի�z(�VԾR��ї�Uz���sUUu����:��U���J�w>ܵba��)B�'�E�K$��cZ. eY)��5˳?e�����Q�f��W{!k۷����n���_#�/o�+���X��T'��1U��Y4��n�ţ�Ԋ7���^��f��3��i&�[�XIQ�ok1��+	<��	@�`�AV7,e�V?�
�+�	N�FM��Gl���
&]&�$�'S󖆵�y�x��(��m���v���r�<u�Uw��h/�0,%�3K�&���&����y|5S]�/�5WTR�p��&�V3�+V����_U~^up�Z�*�@ޗ:�u�N����n�I����P�q�<���:�I�kإ�K<�װI�p�F���%٤�08P[������JX�K<���iF�����	��f\Xs��a\R�L�:M���R�[�ۡ�b����ƕ�LBYVM���M��6;<�u��K	��I��R7�p}�
���ֲU�#%T��(�������
��@����D�3��ĳ���g�׬6��o��<ߐTl�ձ�}:���U�g��{��dZ�ga//"�FY�a/vM����/�t�ڱ����S�������v�T�����^_�~�p��;�㸞;���0����ڰ7n�Nx�%��;��0��{���e�
�y�/:5nݣ|�&L�vs�z�t�U%�)ޣV�8e�Ỏ��Wo�V�)u��j󪼽}���sa�/W|xgF��h���<ʴm}�aIq��$M����[������ȯ�´�&����ǃI|f<?��ϧ��E����R��p��vܐ^Rj�}��K-6y��H��:�*�?�*�E�Y���P��k,�)K^�%c�g�cg'�\]dRO>��J�����⌠p��ݾE'�&�����,�J��?f�^^��$�USE�06��ڣ�^v����}�z7ջv��5٧zw�J%�T��R�w�zuWڻW���a���&M��r���`�FY�W��N��$�#�B�¥,����S�;�.�n�A�G{"�m���Mŋ���"�cɿN��TYO�l(tݕ?J?���e�m��M�_](��$�*��7�m�[!�r�VW� �d-�+-���yT�^�ݿ[���2ۑ~U��n�^A��(2��)��Pi�)n(d�[��gd������
���2~�l�����oi&�2�5�����:��EY�N��䲚R�2��k%�J��ܦ+��%fҵ#�4���l�8G��x4�w������N�����q�>U>�d�m�)7$�c� ���K[&���e+��P�qqG6=`n!?�盜�dlLLd��?`�(ڻ�68����d�M,���`������򯂫�gɹ	'��/�r�l����ݜ�Y�G����F��,���Ŋ@#-��ݍ�*?��3d���;��#�^3>������X��"���g�������M�s�I��x�*�Bs�AD��a�F,9�l|���t�ԟ�&�����Ƿ&��a,��5y%�9|��;K1�.�ݍ�V�Y�!4`�I�����B��J�F_%I%~$P(�JLkz2#:0��\nI�!����v*��R-�+�]��u����r��Ev��4h��V���\�V�f��bd�Rydd;��j���Є�Rh�yK��&k��}�H��ג����<6<�x��1~�}ZI�<�Sxe�b\��}w$�h�e�+#�⿊M�׌ׯ�կ���>�y�����77X,x=�zL��9>��*�M&8.���Á�&���խ�iR���FJ�*5_v���|!բ�3��+��^P�nbd�_���A�đ�TvW=G�����&���&����X�4Q݂��U�����I�)n��W��Q���2~w|��f4W�ɹ��K3J�h�a�,�v�]�VϞ�����q_��e0&e�l�e�Ts(�.��ھ�9{��y�4%�1�<�h��kD~s�1.U*�̣����ӗK��~b�x�a*�u�F��ѽ2dӗ���mz��j�6���.�].�~�ͣ�o�;��j��	q�a���g���Qs��QK��,���8�sU�j^����q	�5|���}�����e�νd��;$�ln/��I�gF��]	*����cUW�*�W>
ퟕ&4���,867)JA�&�Ã&���$�n[y��*������Փ���B��|�IIc@�����~D>�ܜ��H1
��kwk����^Y�\k�ɨ��+n�-&�rFdJ�,k�4��.��w��>�;ח����8jݗ�:7��w�zw�zw�K��U:��I�N���_4X��I����W��@� ���d����
/!r�u��#n�%~�c+'�[~ʡP��C%���Щ+'m�֫z�}J���^�T���gi��Mj%e$-���(e�\8�Zv�?��H>��o{o�e!��ݷ�5�Gi��*v����$8[�I;rT*���le�.���m��µ;*���-ʭ���.�����;K~���j#��FRJ��g�d_-a�M�~d�����K��Su2F��c!wj9{g����4��i!�5��e$H��ϣ���%�ҳ���l��������G+<R���W<��s�+������"%�5��gZ������wrˈ�gvY���<�z脱�����q�
U��ٻ�,�I��$P?z�R}���/�~�s���L�MI/q/|&�\k�Xk�0;5����O(]��ܬ�J�Q����]�o���͕b/��[�6y=5�#��]�`��)�/����0?���Q�RUbA��4iI�h�ՖU��D��������(J�v���c>%*����U�}����"�a#1�ұ�r�h�sߑ]Ռ������ǥ�yc�@�o�oʭI�o�AP+[8͍m"�����3�w�j��u�3]�����q�3I�%�|�2�pZ�誼�V�#�dH^Z��Qc��E�SE<n�m\f�/.�\�6������U�έ�1Շ�Y��.V(�xV�M�X�f�B3V�i܋�Tdd��#μ��q�_M�j`�$\�!����_�^Ǝ�}�v���I���6��Y�Y�ɼ�!;,0#��I�і9��c�kΈ��#�e��ܠ�x5pt<�AQ�a�5��2��	у��<�i����?��|������'ͥ���Մ�H;���\P]w�ʾnQ��.,"�%�T
��qcqwD��~b���\����eP\�]gED�ȭa�s��h�,�sK�K������nOZNkK�/�a(��~�n"t(����^e����	j&���"�i<k�(�W�Z����F_5|�e�Q��k���&M;�պ�{\x��^^���8K�~xW�Wں��Ώ0P7��z�\r���熿Y	cI"�����o�k�dPU����j���z��&M��n��͍}�00?�<��Uy�l'���9�Q<���W���	c�&�D�'5�?��|8�,�������7nJ�SvM|��R��$�	},�b�	rݱ�ۍ�o߯�����m3���M	�����r+���ެl_�OX�XE�>��~�~ɿ7�{��Y�i7��~�њ�Usc���WR����]K��Wp�Z��Լ�K�˥��/F��5gv��)�/_{�[K���0㸴����"Ugٟ�X�z)�wۚ&U'҆��5=�2�����RW�7���ɒ�鲙{�iL��(2;��l��zd?����+aQ��i�R�P��t���)v�����Uj�ݷ�*�+L�x�ڗ���q��t$B�-EB��{�?E3k�é�Yu��r۽��YM�2��S��{����ⰽ��\���w��#���_e�m�v����!%j0b���nB�nS�0�KQ��lr�}�k�����u���*w�UÈ��_%����	YY���5�y���+1]��H�S�R6�)�wm�Dw嗐��J���G�-M�ۋ��vB�x��n.�Ǖ�I�*�*�Q���l���%��gv��ɗ�藗�FwV�Q�����_;��a9ȵlٯU.(���gc�Mb����D,kpԲ7�����۝��۞�+�WQ�������-�W�%�;Ywn�k�i>_�A킧o��E�^�mgf��W��[nX��Q2��p$�(����WnE&���^���K4�
����:��}͢�6VM/&�y��E��|l�9�q�ձ����\_v��欪��_�͹,H���\M.y���D����6>y�׺Ѿ7����/���Ө��'[Mk�p%��^^a������;weQ}��j%��o�j��W���]1ݻ����׭¤�؞�&����D�7U�,�m챶�}���&��I�ll�pH�v�(�yԾO=�b�	������%��^�P���>���ɼ������r�᳂�J��X�E�%����80_��P$��M��{��G��>%i�gc)r).�.��;#uc%�y���+L�M,~i��+m�z2�h"	~G::�Vv��k��r�F_jM�7v�pWP,18�袽w�5ֈ,���7�3N��:6h�1�j�Ό$���w��d�\�n0�����~���J��Q�}��j�W�Z:(��w\=bz�W�0�jw��k�tQ���n溢�^w���y�Ǉ��^�sf�9�s���/a돟ު%�9������]y{�l$�"E�΋]q�/_j�]�ڻG5^�0�U�������}$�#�n�*�Ɨ�W�<~n'j�=tc��<s��cǚծ��a�iuq,���J���F�5�j�.�p�����$���P%&�\U�g8�̏;�xM�3��y7��Z��z�nr�u�)!��ݶ��H�����M%HQ��v�W"�1"�XF�������p$n�"P����R:����Z����d�=g�4�ڜ�T�to�qwU����F�Wo�v�j�ڻ<7��K���y��V_Y|5j��V^��g�^��g�EY{W՗����pջj^��l�Y&ϹB�~�ew唷�����:�����۔7����V^�"/�O�
�u��sO�H�.ҕgۦ�v�wk{8�z��-ZN�t;��ն�J�9����曊۴��)Kn���i�T�l��)do�3�tݴ����A�jc�L�zJ�t��$/k��/m�Gw�
έ;���t՚�_�J��J~�;cn�ҪX�D�M�I)����x�{9Kg!�)�zo*;�M��0얶߿M���65��������U�P��E^�~/�_��+��5JŗeM�u�?~Ȱ��Kс�V
���8S�����*�c��5�tK���Iq�h�����q��XNv�Q���O8��H��ើ�GC���l���f��y�.ۯ��o�s��9ga/��ғ���d�:�J��ո�W�[�nKQ���Ņg+��e��gl��̬4Cv�_���,�S��4��`WӮU�떿*�g����.U�b��6��kvE&�p�\��ul�I�]p�M��9?�2�To��/�pc$����,�hNr�D�qW$9g9e[﹐2��}��\��f�c���XˈZ��q�|�/��ܣ��?UK�j0X2y�V���<����������U��5�y{�'U��5��s���&��/F��������]D���*�b��V��C������߼�,~���"�'��q�2�O4m��o��`�0>�K.Z�����x��^B�(\�mό�ܒ/*KI7T��$��B䰧nBv�`S���_e:�v&�N|n�*���ׂ��qYnX`����d@� �(ν�<Rĺ��y4�
m�3�9��ppv��ōU�g�_n&��n��=����'�95é;PV�y������	�v�������8�e�D��V3���̿�U��袺����O��4f���:�%R��;S����j_5��+��q�â��r�ˮ�W��v�;�qݫ��W�.�W��k_�<�BB@���}��F�������;W`�"bk�$�2Ț�ļ�vE�g�P!)>���WUWڻ�
G�k�z����<z! l0$�6r�|��fa�����7saK݉���qq�6`�2��&<E[��]�:��fo�˭s����&]_��MW��r�Lڴ�e�5e��XhȢV=e�$V��������$Q�z��b'�o6��|����rr��X����"��g&��۰��#!\��]{3�J�Tlc(��:�c����u2s�/G�&�+�oâ^_5[�o�^uqѣj��7�/9�_/;��w�L�����T�vk�LNr�m\y�q�:��~�����ܿ��a��5�Nnq��:#����I,���jl2(	{��w�Ȝ��6�V�yf�?�˟�e݅I[����>vt��&!��Y��l��\�'+��S�E:P�vo�mv�!��U�v�)�u�5;S���{]�>�@�H����p9z�1���²�)����{l�=�nVA��h��6�e��[�W�]��k�ڔ,�T�~w�S��k��6O-ݥp�52|����
E�
��wa��Ņ�6r+���[�e�q۔+%��@��#�,G�{���䭖�)k���x�N�������m�H�hf�Β�Eq�$��z㸂������QU�����j�[�to�*�����XNty� �(u���?�/����m�v����rnY�p�6S{�Xy���ٔ�Y�q.ꝯF����k�ݹ�\������̌�;MQ��V�G�_;&���k�e�d�� �]�) |�`հ��_�O�Oq,��ȖI�4���p6q�p)9�!.$����Ba���"�K�h��vB]��^��u�X�6�>Y�Y_�*�v�>�c�vA�k�;n�h].�����=���F�7X�N�q�̼��_�p�Q*�Z sc��:���tUIs�;��\_vM�siN�i�L�y��_':{	�v?��I����.Y�_o�¢�/'�I����&�Ϗ�Q�wK�U ��o�P��G��4����on�VJ���q���*��\5{,z��+�Q�r-Zu˓��"�B��_[ �%��ə>(ߺn�yK�����/g�.�&����!݁�@����[kR�6�>ts��W�O6���l�����2�{P�e�գ�����Fy������'/Wk�.��U���}$���������V�^�ĺ�jv�㻢�R���v�W�[\���Q��FuK˫�gW������m_F��qݣj��gw�J%��7�ǆիWnݾ�������UEGD��ʪI5��ް1>|�K�z�:<�.<��qkū�訾��XYץ��EV�ըq�j�1�TtZ��E^xח�f�|�U���p=g/V�4Bk�˹��nJ�:�H�ofTb���G�J�9���ݗ�u�ݰ��g��h��]H�p[xȾ�E����/���׫r��
�I��T��e�.B��r���-y++'�Cbwx�6�$ݿ�{5v�9^-NVYX�K�K/���ȳ������/��޼���v��.�|�ݣ��M��xWW��ū\���z�_5Z����F���m]���6�ѵu2d��to�/F��e��Ѵ���s	/V�;��.�K����_g��c&�4}���ۧZ�bf��Y���ʨR{��N��rϲ&������4o�L�>L��m�ʬb��p���J?�M�\�ڙ;K~B��u�K�"҆�����-�O����(WʡQ�C{N�l7"���n�B�S�l�������"���O~���Ն����H�<�nh���	g��D�V/�X��P2����7%���"��D�%oiZ�UK;��Cd-��V ����;�f�*B��nܿ)��}�J�I��n�B�	�/�%����/E}�%���&���5�-{l�/&�Wɔ�l^/��l�ä��4�7o�x.�k�0�@�뢯�������y�\0�R������/�<�������㺺��]D�UVkUQ�P^g"�`�U��nʹ�?,�oܕb%�X݌��۱�J,��탊�Þ��Q���V|l��!H6�UIk�3�̈��6�=���p��%��2*If�|*R�䵺�޲Jυq@���`X�jɼ�Ŀ˱��g�]��z⫬��W�R�tI���dё����6{�Dn�[�Ly�Q���D��.��C�=m(���oc�������S.�K���K�tK���Z����I�j�j:,~�Y�a��qqW�9��Xl�B�]݂��`�I���ёD�n���w�Y*��"��sN]��&��*����P��vy-[n��4q���H;�9,~�0w1z�o?uk��RFm��ܬ�~Y�5y$���4_�=*�@ψl�y�&lK�X��nzYj�'K�mȓjbx�J� �-�g���;�6<��uۖ �e^��\;H����o�-i}����&�����X�|�Y�ׄ����/ck��_��04XL%S	��aQ����8,�i�&�2Y�&�_��[�.����:�tQ���v�W�[��ѵz�yz���諏EZ6��^k��\ty���΋�o^�^w����ڻF�۸o�^s�QN�D����9���ﵣ>��vv�ߎ���޷ڻ/�o:K���q�U]�Et�q���"E�
�5S&��$lN�=h�����U���5[����v�kY�n%�3_k
��\�|���g�|���{T�h����	�_E꪿p㳄��c�&�g��?�K�ݖy��"�Ł	
����2�zvzU��r/��IQ��"�O��~Bp��HY.�\�ٹ�E�"�vV�T�n|�M��b�����2���r�K���1�UU�/uF�����V
�����k�\���z�_5Y|�e�U��V�:5qѣj�Wh�G69~z-\s�ן�=~�u���]}[��Z�/q���Z0�L&^��v:m����ҳ��t�|;t�Go�&�k��R|��l�ę/����'���_��ò��#r�"҆��G���:Y��]�ƛv!(g�ӿ�k��,���vo�4�-�p�p4�R}X�%n/���$?��nw����[v���W7-����	*&�o#����e�q[tA`ㄳ��«���_;,�`\�f�M�N݅d��PۊM,^[aN�l���KW�/ �+r����V1}�Z�(�����I��s�y��6�BA۲�s�y]-N�'%��GkU�`��a��|d�o�1?�)"g���:HJ��~|���$�ľn���<��Y���������Z���X���qk��]^c�a��.����k�'f=|�N�YT�΍|�[�7�c���h�Ϫ2���;\Rf�����Am2X鰨L]R�ֿ6˺��2T^���=Z���'��tO>r�4��nU۷"�vX�ʲ7�i��+�L�i�[�oY<e&|�Uۻ"��\UQ4]���*%��SE[��Q��w��?n,4��,�mO�j��tY�Xrj���RZ��h�q��e�j,3c����<~n.!<ݣzl=q�QUU營޵tK��㢗�o��%��b|�����dm��YWD�j���_��{��,��X��Vq�-_a�&�*ے���X��/I�F�KY�_"�Ȼ'�"�qK�F��~�>�߯�z2R�j3E_2��zڳ�ßIIN۱��;,R}d�����M�|�2��e�噰1w-|�lM���݄��C�ʨ{�w�@�n��_qr�RK�n����"A3���M���_gp���u�ȯ�j�`ZK0ݑh@��|޴�E�q_�7D���걔L*�e��Zf���y���k�;����UD�](�W㾯:�������v�t�˨˯����7�/;�o���(0P8tK�_/;��w�p�w�Q.�S�Q/_vr�jիT_}��hǚ��WUIy�O�]q��D��	qaw�]����{�%ğYag_/��覻j_����n0���2W�w�d�R�S*���5\֒�S(�z�r���Q9���g�(G�k��y?�x�
)~�j�]����5��:��8�F��
��2�h�����(�����#�F�Õ��S]�bi�V���L�*V�S6�|�~+HU��9�F���s��矁<	=�&�����m�j�uȑh��0�U�yy/v�5o�V֌wz�����Uu|���U�����U\tj�/�������F���p�W5�����я�Ə0<����	��f�~��˶�M��YݦO���v����H���kx�E7M��[>�v�?��a��φ���aR�#�P�ߔ0nR����0��ly:�\��iQ����U��zՊՏ[VjK�M.����%KVT�dݕ����*P���GM*߲�ȷ��6��e
L�T*
MɎ3J7"N�j2��v�7i�ɒ���ƕN�VklL���r�ܷ�C��r}�����-"݋�Y�ʷ)�;��6�~(we���I�A�nD$�)7&h�W�����,���ȵ�9>$*�%dn�;8i�-(l�n�p=C���<Gv;	"�H:��.89��a���ٴ��JR���<3�TL$�o������%/uEj�$��6Mcqqk���8(��6r)d�O'����ғ����w�'_?�-sÛΏ���n(��;���u�ݐ�p�������"џ"���i4Չ>����V�R���$M��V�_�n��e�(�E7od�R�I�����6�Om�R\cҖy׳�3�Ğ�7E"����܉��BI�+�p4��p.Z�m|>�L����*����Uj&�3Ǭd�xo����r���4�0�U]a�qW��'�)
?�(V0�@���z]j5��U��tj�㗁�<<�}���j^_Y|�gUw�z�����D�Ŭ����ά;�UK������.����f���	�������W;��|�X`�.Xr �;,."sy�j�ˬ��V�(*uw���m�ы�5`�+�����>�4%�32�<FJٴ���Y�<��c����V,�.���4�|o���B��Cn����-m;a"��o/�����~`�-�<�u}��X���{.݆���5��4l0�τI��ȁ�r�������BEq�b�Q�c}��e[��s\X�Q���m��nK"t� l�*�cZ--}�G�Z<���V�:7e�΍�ջv^����������W7[R��Î�wj�+�Wn������7�/:6���/k�6���������o�^s�]/(���ꗮѿ�yyyy�s���n�ǅt���^��u��R�y/=��ͣ�=���+]q�}��
&�2�z8��9z:<��q/��'��=�\֗��*��q��U[הf����I�&\a\K�]��D�\�R�h+U�~�Q*�jl-=_e�8`x����ȼ��)�x�ƕ��%��[�Gn�;"�����l����{��3�_@�\\s���ſ�V�@�K7�,n[v;�X�R�{����N��JW-4��N��¹"r,��UQ����WkXsZ�ן���u�w���F����|���F�ڸ��櫇D��qѻ���旜��~�mK��Ç9|�%�h���_�?i0$�7-��\�%|��fRR�e,��fΙ �C�u�#�1Z�;�"��^)#뜥VR��-y+s�^�R��=�R��W�ǁ����-���bd�vJ�Ewk�r��r��[?9m�+��L�:��(�*�!kp$��l������g��[r����(u�o��F��+|�f�;d�&�'�Ȉl��h�-$v��_v?��V����n��M�M�\�vQy�nY�Xݠb.U�d��P�S�4�fN)os�qxt�;�a��^MW����68I_�}n褳υm;�������Ku�+[��V2[(L��:����c�U���q��W�m_b���Oa���_���v�\\c�yz��uǛ�;\���/�4�lu�y�``D�AB}�qךly�s�ѣ�8H؟10W���2664���6#M��a����6�����d�-M� �V�^���V9g�(�*�x(N�:�<�����s#�������V�/F�"X�K�j2��E���'�I�$�|�.ș5|gޱ�\��c������0RjL̉d�����5����f�V�y��=p��q�̈́�U]U��Y�z7�{>x5c.XTyո��7��ʬ���X�(��x�H�|5e���;Tshâ5�tWJ�j5���a�q�ۊ���>�ۇ[N�Y��
�"��9T=��˺ݟYy�/���h?�	ہ�%P:ȡ1�Ï���齶5���S�T?wg��Ajb���vMŁ&ϓRY�����f��Λ�<���_�Op����^���&dMU%�e�U��Q�����I��=,V:���d��,��y�cnYh��/"ۯ@�S�����r�_'�F��F�۸7�����Y��B9��@�y�Ռ�"���4}&i<ş�x�p! p~���ѻ�_�
��m@��ם�z)�z�4jݾ^uqݾ]|�_5|�j㻎�
��R����uj��Z�>r��n������������^w��uJ%��o�j�ꗓ]�x��eٯ/c�3�����sK��WD�8�V7z�s����y{G�xn-/O��UF��\h�q��5j浇�dɯ�V�<=~����I�X=�V6r�I��2U����Ɏ&��5�\�(�1�XKE�UK��p���"��N���`�F�Ñ�
���b�z��+�sU%E��R������ky}������r���`Ci��x�������)e��&Ż����t�i/I߉����*����"�Kݻ�
��Q�to^�����V�y������Q_/<:%�ᾍ������/�D�\tn�uUqѫ��j�����/kF;Y�K��v_6�,8���汓g�4��&�;r����d8VK/�N�ϧ`���1r}̗e�{�[�B�R5�O�e�����wd9n�x4�?Y�q�;fq����DVR�[9Q�\�s�T�5;{�����,�r�v��0b�o�4��c�)Y�2��(��J��Ҭlbwl�s����Ѣ΁�m��k�W�L��W,_��׬m7$��c��!l����7e��W�S�\�ZM(��&/�B����.�>)g�d�z�NW�n��\T�d�r?�kq�`�Rik�HKQ:[u�Ⴕ�Y�Oa*�J����Dd��%k0._��nW&W+	�����FDNF��J��$�ݫyD�V��7e�ݣj�\tn:��	׭�:7�<x:�P��6�c�q������^wջq笾��sc�v�qp��֋PPT���n�>��4�&U�������`BBG����"+lnD�L
����i��8m�t^��{i�|F�S,���q�FpQ��\\Q�Q�o��Ϝ=t���n���n�H��~��	,�I���5��-�:���a�__�_"�K/���//_�_�|L�Wz*��].s����f��@�ί�R�p����s�WD��?:#%���bo�;�r�ᗿi|:%�K��a����j���<��s���|L%��(�e��Z�o�1���]n��W�U����u̸nl�yZ��'�E|ԗs�ܖI���^�K?�e�X�H���DA�w^�I��Nl�MZĕM���u�Fï��b�����o��X�gX��V���X0��� ��a�؆~/s6T�p;x�)]Cd�����^��<�1�	UYf�e�C�ԫ˖"/�U�^M�^MΓ~M�X����|e�L�L����[�rI�I�n��FfFZAUD�B*�h�ұ�,��U.�@悱�]��ϝ[�ѣE5���V_5Z5g}��)|7o��Vy���q����y����5�+�Wh����w�zw�zw�z����]��D���Q]�}�jիV�[V��7�j��EW���`b|ḵ<7��/G5[����Ek�=�ḵ��?�0\�.�_��i�Ѱ�K1�曟����&�j^�5To�������}(+ߴ����01�y��/�2�'6k��WK�P9�J*9����\_�&ܔ!�=���2x��AI�rM�)[y3�XM���nJ!��XH\H�5��+io��[��w;m��u���J�X���ϗ�X%Q7�X��_��ēF�� ���Y���W������^�5jڗ�j^��e��V��+�Wh��]��Ev���_uF���ݵ���v�:����-a9��q	���=.[}��l��O/�&�k>�^����|Q|샬��d����v6��>*n�;����o���ar�ȶ�rb���v7h�7S!岛Yd+��)HҪƷrP�dS��xV��Y��d|����~Vͅ�����*�����n�[�lm�LwJ��Ϭoc�o-Z��e�]��#�Lߒ�hn�ݝ�T���ܕY�w�v���!e���in۔=��]�\U�mN�1����O+)l��rr}�l�nB���tI�$[rM�ݏ�xd-����k��ݶ]�cM���mE�e#n��ۖ��P�����7" ��_�AK3}���c��b�.]�s�lv���͔��}��
��j_�i}q诉���	T�u�4�n��u��ͅ|llL<֕h���]mKڸ�VԼ��q���VԽ�e�h��&�dno�k��������66lh����Ȗf�J�9���v����K�E}�m@�,{-�ڱ��2�)#$����_JN��V#-���ݫ��n����Ni��ݻv��b�M��,_����tqo�qvܡ#?��Fj3_2�/9ڻ~:7㢽c*�B��z�\
vvR�KrGYUz�E'��*��W���:�q�U_j�t�5[�pի/F�[��ݵ������	p���C�bz诂��Rf������nr�SZ �:�БP5�쿎f����qI��\����F�*�JW.v܍�UnYm�D�AZ�_q�"������׉�a
���v^O���|~�_�*�IU��ye�?����UbaY���[�l��|��^���g&"�MjMr��T}��v�=[�_^�j�n��H<P]�$���]uBo�|�p2��7�Ѹ���,�}$��>vw��3m^�|���p݉�vÚǚ�O$�Y�X�Ⱥ�AU���h\W��_�t�0��F����5�7��/�D�Y{�y4�&�Eq����/0��9��k�5gF��՝�+�Wh����Yѫ:5gF��՝��Vtj��y�/;��|��Ѿ��ݻv��8p���΍�L7���U�tp�Z���U�tR�^����6
�&�\wڻ���o:*�Q��kW᫏�8��W]�.�z�e�W?�A\By�j_G���Z����ڪ�G�$&h�<�! �ԉr��<*%��^x�`P2��q�cVE	k>3�܉�i<
�G=Yd��
ÃIG'e%nF�"mhғ�~[:v�g"���2Y-������[v{M�쥃���ݰX˥^T��y�D6�ʥ�K���{֪�.�to��F�ѽvk�h��]��Ev���+�S�}����v�:��a�q��;�<�(�u�q֬?>sy����J�i�\�&���ۆ�mӥ�<0�Ƨ��	'�p�y\��N�C%��!J��.�!l�k�I=�
M������@��,�$�N�ѹ[��nI_�U2E�iS��9\�ϻ�����a��"ˑN��[}(V�J�ä/E���oe�V�����/�����:Va�<VG�~<~�?���q_N&����Z��ǸL{��TqX���,��rd�T�J�N�Ct�xVWѥ�Xn�3�T���[r՚n�H҆�t������������J[	iZ�\�V<_��!%T2.�j�*��@��©�q|^~�^���'�V�~�[�S)Vݧv]q����)<�%r��w!.#!4By���m��}��	����xtK���O��p�q��}�X�J���ǅ2dӣ|��߆^�;_�#eZ������+���
���4.��3�sE}����Aỻ`�@��X��	׆?���N�b�_^E���ٯ�����ٹŻ*��������۷n�F��oNk��D	ݺn|�X6z������r���=�XK����߆��������7�y�����J��V�^J��v�j1�,w�]](�@��j�e����/;WUoQ���gF��L�E'����K�s�&���jir���9{�ڿ���;����4�'J��5q�s�j_�5��7nE�(rZ�qDڋ��S�X?���%Q��J/���#.Rd"�l�N|�7��=dPLiT���� {$�<9���J۷}'4�yRc���J����������5mK0��S�[K�1�[d_�qw$jE���m�dfX/;�ˍ�H���5�g��I�ь��s!&�3.�_f0���j���pa9�Aa���_�.�K�F&Β�:�`�`�>��F��w����j� sh��k��o��2k�V���q���=����Fꬽ��hջF�۴o�F��o�F�6���՗�V��5nѫv��Ѿ_5Y|�j�w�h�}��s���*����^����:3�z��j�y�/K�����\j%�9��͆��[R�mK�V��d�ջ/�[R�mK��V֌pQ�4��9�4&��5Ǟ�y���O*�����	����������^�2k���gVԺ��j�|MX.w`�\J�z�XF�i<��M)J�a>˩:�Y�ee���HJ��zRh�m|+~ηm���y��~���ϲ�Ɲ���gp�}}�V�X�+�8tW�N���TWh��]��Ev�uJ+��������޾�Y��k\�0��k�[V���Ƌ�.�h�qq���O�V~�%|����6�M�aك���qm��+{�M����z�����I�b��;����O���uv�~s�P�ݧR`�y+-�o�f����_���������H^�̖&�������M�+�R��$mʛ��d���N�����ov��[�-�����~U?DVK�|h1L�x��d��|xԭ���~�[�k$��w)���i8�y��6�7Y��k��Ie�X�y��@Ȩ��f�܄�E����T��ݭ��w1u�r��/a(z+��Tv�e���ӵ�Jnʟɋ�k��R}�^9f��(�&m~�ˬ��kQIcL���<����{(H��e���E�׬�srq֒�i~wy�ǚ'��(O�Q?�~�K�¢U�j�E�h��<��������K�z�Wq���qj�<4sc�������B�!Q}�������Բ���PZ�6�a[�1���N׌gؼյc��jw???"��-�	4�2��##o��r�⍤���Ti޻�����ݾ�ׁ�ϟ??�y�h����<6���X旫��5hݗ�VԼ��x����d�y�^Z��&q�Uù��b>��.�R�n�Q}�����{�3Q���MW|�q�椑X����4�V;����5Ļ��8��i��]v�EU�Tb���6
E�3����l�U����aW��#���P.��BqI�kr}�>�������f��_��O��r���/���q}�vJ�\*����E�&���,�ۓ��Xu�Y�܍�*�9ff7暁O��K>T]
�o�2�)+�����N)>mX�Z�u���&�������/,�������a1��e�ɮ4K9���6c�۲�:5�e�?��єz��vYxs�%�\�,0��y5�]��x����5n�Q�w�~~t@����7\xmQ�/|��j�w�_5�Q���;�o�F��o���;��w�{�|6���գV��7�vs���:4m]�����v�� ��qѸ���	��xo���:3�|�<7ں�������Uy{Ũ��϶0V��^^�j^toL�֌tpջ/E55`a<��}[�e���yM'��F��.���3������;Ugj�$lM��
�o�Uv|�����c����Nz+���cy%T����n�܋A�ܓ,y�oʿ�٩4[�g�&�o��"��H6t�D�N��5k-�R��[b
HF4�#?����0e�0_�9��dNO�Ύ�8����Tpڣk�Xn��/��\tj�}��W�_u}��W�_u}��Tjά��mQǚ_6�:.0�qV�^tn3U������6�Z�4�|w��$Z\P۔C�
��ϋ仲��-��7K�P���4W���,�k�|;q}6e�>�M�ld����ל
Im����m�ݍ��w_�[�m�Z���=�̳�^����=��i���������Hە��'e63J����*�'���Vt��v�����YHw��Ը����ZB��yz�1ݷR��l��������VR?�����5+���;�r8�mʿ,�4��O����m�;�M��_D��M���vV6t���g-�V6vR�����Tψ�ZH�k)���O����9]EO~B��[u�������o��1;�d1���4��M����FF�c2|�c�/W�����@����\tgjk��3��4ߴ��Uo�j�<r��@���F���>������^wsa�־���e,���*�X݋�|��K�����Q��?��Y������]�dK��`PP;���mc���H�0t\u..5u����n��<ք��&Nr�˩�L��F�Y�n�n�L�w��:��b~�Q%�<ֹ��h��^tq᜽�
L�7�4&^���g����x>evX���.������<2��������ݾ������艁��E9���h�����6��E���aU(��w�%�X�5n%�΍�%�<L�Ś����,��Մ÷ոYڤ��Y�n^nR�{��e��µ��`��*v��7�͢��<�����-�#KY[���cҍ�פ�����
�K2_�̬B����1��H�D�dM$*�^E���v�U(o�⤞�L�+��f���>&2�&�vM�a��%zOu��D6��:EV�X)t�f���U�\F�K!5�0��UP7����?���qea�����U&��ܥ(�V�f61��O	�B���|�n㢗�����Î5��z sa�/F��|�hڻv�2i޾�Y���N�dɓ&�/F�[�h�}٦L�2�D�Q_vs�9�s�>|�ի}[��1ḵ;WR��%�u�<7���v�WR��qk��<*�9��R}������f�4�����H��sZ�ǆ_ɓ]���5�ɓy��z�Ea�t�U�]zy�ځ�9z8�����li��D�YȘh��wn��	�'сFM�Mm�U�FFC{%R*~U�U���/�%Cm��Ym�ßI'�p¾Z�n�_e���H]y5��$&4Nh(���P�i��4�U�&|g��])5�W��w5Y~xmc���Xnᗾ����n��F_5[����������Q�:���F�:��K�чϜ�08�.0��W6:�9ځ���'��--ͻ<�*��U��M�H9o�~J�ܫ�z�f|_n��҅ed���J��V!�܆魲W��֓v!ku�e*=l��h�LR���g�b����d*�;=Z���T����:̧�YX�H����n�o^?ʓܱx;�Uğ�/I�N�,�b66�\v��l�[Ze����j�N��E��y+N��3��;#d��+�oېv}���$��ۭ�;d-�|*R׈J<���{�ro+��^�Cg�bm�;�_�zo*;�e08q�TwcL��[���e+r����������+m�R�DW�J������R��T��Sr�j?2��U�km�ҫ���7_i�Œ���c��,��ߠHY��:��k�ٔK���<<�n �#+�α0�!.4B\s����G?9��͛��0]`c y�\K��<2��?ʷ7m��
�X�S��+^�g�V&	���#2$�wsnK4P5h�J��ʒh&�5n9��������w�ɾ�Anܷ7w;-c�.ժL��Rs�\�L��v�7o�F�[V�aÄ _vw���j���Ɗ��N^��[R�mK��i2e媴�2~J�JE��?0P62�IV�g&���Xf���}����/��<)y��/=UL�\�֯a��mc�q/�3뤼�s�q��M��j+�_����a\D���B�/a���\��EUau|dm�䪭�;�1�ȍRfҒ�Y��+<���u���x�krMN���JP��"6?���q�a(V�t�f�#Y��[d\���e��mڅK*�Fc�F�ݍ�����nn*��>�U	w>����7I���Eƕ'\���jȿ�P3Ҭָc.(�w�R����Z>����ׂY�������	�ڵaq���&��T���_��Iv�C���}�����0�n):���\Fs��y�旚^iy�j��tKѵvuS��j�mn:��iz5f�w�zw�&L�5�g}���dɓ&Q(�J+��������|��s^��68ʥ�ڻ}��sU^^](�R����sU�qj�\r����F�Wo�v֌x��Ú�5gF�ɧF����D��/E6֭hƽ��^q�o�.�V_�Vl5|�irqRH��ʷs@�y�����6hO�>�&�qΌ6j2���K �dF�ȍǫa���Ӳ{,o1.�g�ѥ%D)"��aYύ���c�k�b�h�6�0)�	<7m���9}�SJ�K-!D�nP\:�u����c���U�7p��V���ޝU�7�j��+�Wh��]��Ev���+�Tjά���n�F�:��ո�i{Xn�ỏ5�|�f�ч��(�<�J�>��O����*��;,L*R��v4�ƚF��[J޶�X�q[u��wj�ȝĉ���Ċ�"�r��#�m��*E�N�r����*��v�V|Tݻn����B�V���)�J�I[	+aQ��jp�_�J�ҫyjg�����?*��[!�T�~嗻
��k��l����e�w���YyT�޲�����:޲��N���Ȇ��p����X��Y��ۦ���ܭ�$��7M,�҅gl��~�H�r�1M�nǊ۱��)+�S�d���v?���V�[��c$mw��v/�Aܐ���T���T���t���~i���.�^��קwy,�{�;��M׈l�ފBP���n�캟n�g����]��xo��^�k�tK�����[���d�y<M$g8K���|�@��'>���誢��G����j^xe��D�vk¬�_�)4��|6/q_`���3s�����6�bE�,��YW��y��?��2�����O�w//.ݻ;�Wh��N�\wΩ2dɓ&��F��nݻv�[�mKջ}�f�2e��^��R�ѿ6�xmK��W<֠y���3�%��yߎ�w�k� �"e�-_��\���|�a��E�q��Nz�F�f��a��yT�]%�D��xe�U���\�����\��֎�,�tQ�5�5����a�݌����	�8Dg�+Sm�ұ��%	G�O���xv6Xn��[ቹ`F�.J��Un�B���E���r ��X�26�M(rO�7_�䍫�]���_���cWGl���=��h�n����;/%�;���'X澾㭟�L��2:5�z�XXSt�c�u��.$�o���WḠ`u��Q䰄�i0z�����Fh�U��FKѓuXfD���:��;���&�����ȮX(��M�&�,��̾o��y�/��j�^��jݵ.�uy5�n����X=ts�F���jݻF��o�F��������zw�zw�zw�zw�z_5Z��ѵv��ջv���|�0N^�]�sU����uy/5���zxo^^K�/5����y��2kZ1ݗ�:7�F��D���`I�$]���cc/��o����0���uZ�W��wV�Ej�h�sc���G�D�Z��l0=sD�3Q��̪�&�*���k��P;�:�jĥ���Y(������%~]҄��D#�6��+0�SV6��}�������� �|�g���f��ù���@�AhƪQU�/F��v�㗿�ӽ:��o�����Vtj΍Yѫ:5gF��՝�+�Tjά���n�G�6����5�z7ݝ5n ```���Gk�4j��H9m�����<�������M�������n#Q����ې��e.�J���!v~J]����J��v
Or���:�H���ҭ�J�%be-�v)��i�L�-����VXM(��7iI�e�v�d�v��p�X��v+��Ǭ���+%��e�z+�����&�(e�u��N�Ң�l�J�����7v�M�ֻ!��T�������=�+�e�Cr��J޷̋�#�J܏�t�Y]��Ɓ!|�-�M^�D$�������h�q(m-��.(��r?�݋��3��MoYO��)���3[$mw��6}i(|�z���������7����6�z�Ⱦ϶���{b�[��L���vK�"�^Y
μ�Aj©���wє�߅-ZM}�����_6�0=s@��qkgX����5q��q��'>�s}���������J*����/��3h����ϗ��K;;e,���c6fvщ�j�2�i	j�f��

&6��Ytɗo^�/F�<5h��͎�%�yyyyrd�Z7p�:��dɓ'5�j՗���� �/F��L�2�۶��&�M;����X�ɳ��d�k��Q}����UW�;�˥����f��E��W��Ն����ḵ/��j�m]�^uq�ͣ�v�c�F�����	U>tj��=US�v^���ޢ@��@ɡ��*t�Ej��2�Hn���[߄�FXqH�ɼ�E��4t�k\j���Փ�n���D�j�ۯ���XB�g,�c�H��.ѠI�q��L��(��������{��k{�d�Ԫ����7�rY�弽]�2��;�2�L2���`���FvȺ�Ʃ*��ю�3�9���J��=��V��v����~�ly��~k�)�:�i���&:����}҈j�k���h��Y�kס*㰸�'����l���g�W(��G8��^���/_V�5e�ի/F�۷ݜ��p՗�V���o�v�[�ջ;˳���F��o���5n�V�?:4@��qk�z8j΍�U�/VԺe��Xo^^U.�Uq�K�yU|�ח�Wpޗ��T��z8j��R~P!X::󯳓W�ɬ$R�Ie�H�z恸�I&���I	W���|O���O�?`mFBQ����3D��%�Q��2&�^s皯���y�����~��a�Բ
s'�!�aq*�v��j���ϱ���pq|=�h��Gn~ʚ�f�iCr{	B?�>E�"Ec���*By\ch��Fu쳗�D���GD%����kFi|�n�՜�Y�ệD�;�Ue�/}Y{���V^���՗����h��Q�:��՗�_�6��G�Ɗ��W���	I'������I'���ؽgw�?!vE�-z/���e�A`p��yR~��h�[���q��m{n�C+�Y�X�|���E�m��6��l��?�Pנk;d��+-� �d���T�����h��F��$j�K���$8nʵ���k{�|_YZ���^ѫ�j�����$���Wa��� �e�/vߴ�|e���'�wj{L�{g���net���?�M�[�콖��o�!�;+v�7��[�a�'�9$E&���ÇJ�܏젥T�C�����I�����bc���fB�[�+{�I*UÈ��J�;V!���YNK.^��o�2�q}���ܐ��V]��CeN�e8�����!���E�ԜT�ĲU���Z�NN�@�r�k�/�����h�/.�U���o�v��9ɬl<�����z*��Ѣ������s��	ή��㣇�j��U�'���D��jd����86�!h���^���Lrh�2�8דK�˧;�j�͎�;Kɥ�ႉ�aI���I��Z�j�	�M}�z�gv���}�o�9Ϟ�� �v�۷BdӼ�5ٮ�vk�9���ͣ��MkF8���5��oK?�W�g���j�n-c��r�3^]0ѣ�^x���w�l�]^��T��w�c�k[�S�/���?�;��/��Y�f��w�O���^�D���W��t���W(�5��Q�)6�v��g��[w.�F����O*���;�/�O�j���|��@�Se,�VO����]?S!kɹP�]��ʆ$9���e�#SA�H��1-d^�n~����@�ό��������f�}�����֊
ǜ'��>�I��\�%�_��Cq���FY�6�;��/Vtj�{4&���k�Y���u�I������B����V�`�ȡ(���c�;�����e��/4��/j��vwh�ѽ5�n��B����
d�٠n%��L��5q�����Wqў�Kˮ~tF�).�ѫ�_ū���j��tR�^]�d�sZͣ��v��sZ���N��z7ݝ�z8mK����FF|���>U��<�7m_��y��_�����"����Fj��	����3?Yq'���X�Y����h�ɫॖ��f���Q�漫;�tK�u��o��\�ѯ����������ʤ�i `pln0lcx�\�$�,��)S�k�)5d�����l�\�Y�� ��V�Q���?�����f��//qj�WgUv�^����k�v���W6:��g�^�v���v���Q�\�0^z�c��q���a:��y��j���9����Fs��_�XH�>f�B���+�6�*2E��r�vD6Ზe�n&O������FK7�?2Z\��fBY�M�jnU��DC;g�%qH;�c!�IT�n�+��C*g����v�*�*�^?����lN���eq2D;8��[;#C�{ej=�����T���l��FN˽�eu=�R)��y-�*;�aes�⿼�j �R6�o��Et�xv/[S�ei���n�[
�S5���gn"��צ��k~�����\e�P�䔤_�-6&�)wm��'r����[aR��Y��l䊗*����5ky�-^I+4N��;[���.R^/���Q�uc{Q�z*1dw%��␷#�e#5�"L:#$�*nW�!D$�o�W%_������$l���ڟ<s�/;�/V��8�H�y��c��F<��j�ix<��Z燬%�޸�sQ�V�WX�֨��I��[��=k�`l)3D�O�=�tX������f���/q��yѽyvwպ�4ɮ��Ú�lC�so�kR�}-����R뷯�a��ī??5Ɓ}[��u2e��vi�&��9�ѣ//////F��`F�x��ѣ�^�~���I�]��>�(�e�?�m\hU���d>��ڗ���&��FX���q筯�e���q΍�n|������vԽ[R���Ωz�y��q��]��qݫ���W�P��{�3��Y�W�*����	.̻.������FUX���Ґ�c(�	<�ÛnL��n�T���|D~���X��۳�°u�z��������[ݟ%nD�eR���^&�b(�~ϟ��˿!o�������_���ֶZ�)c���vI�x+W,��)V=y�,�eR�2jId+�O@ߟ�&�}��B�
Rזm!W,Z*8ly���/���]�������Rz08Wo�i̗c���� ���ÑG^6�nEIۑ_�,�,�V�^��P1�|����l7��&_zs��7j��F���˳��֏=e�cQ�y2i}���~�sZ���xq��΋�讗J%�^tsU^^^].����s�v��ջV^�iޫ/G�tӽF���ݝ�S^U�~�y�:�]�e�tU�q�"݈v��;i%Vr����qqI/�E�OY=&��x/6�! �Ry7f�8�)��/����Xh���͌b�[�ڿ��9vj,�h�s�"����X��������gc?����`dT�a:��XiD8d�.�r+<*/;��HN̉��n�8߭��>x��@����&�uºa��]QZ�i|v�ᗿ����V����ݵ��{�a��4�[�}n1��w��>`t\s��7�<�ڣ	q		�27�|�O	/�4%��vE�
�j¶���d6�Y=��K���}��B}n汁����y"���IB�V��_��۲��%,�De�N��51�ܬ��%S,�ڞƟR�Hu-�2�M�d�?%X�Gl���I�l����C;
��v�o7�����t�^�Q��d>KaM���[~��s��)�{v]�w+;��ou��������w+<�W*� �$-�W���56�n�;Z���i#�J�ë0���dS�pݕ+�J��^��;��ᒶyH~&��ۧknU��n�"����ەo{"�J]ejۋ�Y��8c�M_̴_#qS{�)K/M���DRP�ã�V�#ۈ�ӵ8��y��%�c��J���+�OՋ�)��n&[�܈Q��g�109�:ፄ��3�8Hxp?z���FX���V�Y՗���;��D�?:9�ц���to�v�tTg�7��	e�|n���!*��a�k��sD�K��W��xwy�a�}[��ӣz�e���k?w^�X��Z��=����wJ庽W5�[�y椖W�vj�vj��F&]�d˳���&MyyV��5j�V�۷�����Ϝ$$'^�q��k6m`Uo�E�xy���&������vtpջ/F��~w%�ջ4�<*7W�.�w6��ڸњ�5�z2����F_���덅��_��UW�Z:%���,��q�z2E'��X�EY~�y�\K��y��\#/�#����=ܬ7�ie��gѕAK)���eS��k>1'���,�S;�����ۖ"/�"�����ɩP�D�K�V����nG'�ˇ~����{���S�=�(�kgj�*qF��Cr^�T��e��Sd�*�n�Z��j���V^̴�߻�f�WڕH�a�wK�~0��F�	�A���o����B+迮�Q�֌�Nx���̲'̊7�"������h�3Aa����\�PZ���_tg��Ϥ����������'�a.�����6
���e��2e��W�2��\�.0�Z��S�}���Q�V��|7�y�G5[�]��׬%�WW�W��t�����/���xn���u�I��E�hջ/���hջ/���y�Ѿ�����&�V�kʷnѣF�۴e��!?��$�8�f��
�3Dd���y�q��l8�,p_�̵V|��������F}����EFs�V�l3�UV�媹����������q�ۏ�!%��`��d֣!K���WK�uc!0��:�UK�)<��ʣ�zt6U"h«{��- ma��/�ut�a�E:��R�g/Vr�g�^�2�ᗾ�{�a�k�2���wFi~����/Vy���q�Fi~������f�F�OI*����59~�78iݶܯgm�N�v�4�-z�m��X.a���g*ܧ~V55���B��+�γQ���5��Q�M��nHT��-��O�R��[8��' ��V��nv�I;YV���˳�婔�L��)l%T��ciN�ۿ2X�fN���,�JV���ߔ=����-��|���E䭅�/���q�r�jt��R��*B�Ge-���N���v6ܶR�ʎ���M�>����i�U;cn�ߒ�d�+k�z%���/��{c0"\��$7��r�;?2��j�58�W�m_���{#l�Y�V]]�J��~Y}��C�w�R��cc�e�nJ*v�ݕ�T�_m;-��䵸;�ؚ�s6nB��56��i��m5��~R���������&���i"|�X������$g�<	dm$;�p�``|�ǚ_�'Z6���/��ծxh�}��ڻ~:*3����n*����̼5[��юD�_�ځ�j��o�/Fw�/&MG^p7[���:l�!n�\�浹��)e��;~b~��j^2���E,��ב`٦^L�z��y2k��7�V�ڷnѾ�(ѣ}��s�V���WѢ///N^��'��=�$lM�����qv^�i|xq��F��ѽv�˷�њ�<j�o�W^i��ї熮�z�%��Z������Vיu�[���p��/����{�#>�F�����㤳�����hω��,��ɢ��d�o��VM�͹����_�����Q��uF���_�)E�!��5���K���o����H��?-#P}�}�^Ν����3�ߍ
;�62W~���i��Ȩ���J\YyB&J��ձ��Sm�|ݺ�ϑg�d-�6/���"���K�) �s�ʤ���3^^�c)d5m]��I�ѓK�|��o����M�>��E&9g�;�s�0��a%�	F��{���ʾ�%ЗsK:��}���8+7|�Qu�����l�N����������V�d�֠y�љz�W|��	k�<p9��/�����V�j�y�j�]�)�
�'Dk�o^Q_/5�uk���?���_5\:%�#?�}��5���w�ջV^��7���^wh�}��vi�Ѿ�<4jݼ������Nusc����I/����
�W������`H��İտE�{�֠y��i/u/v�kY�ng��e�]���5�R���q��kI{�����A��W�K,$��0��UTf�E�^���|�/.�W`���D�.��ʤ���,\����.��j�ۉxNlwUL7��V�:7�_u/Vxe��j�����a�Z,2���v��e﵆���n1��͎��v�?�y����L���?�u��I_c���,����7�n��n����$d�r���N݅d�%�����Xbp��H�b�5�f��S�ÒՅgy+{ݔ��쥸n"H���X�D��M��P2��io��2�}�,N}
U��\y�niv�P�_v����Z�o;��B����/w%���2pN^�M�ֹ$GogX�V�U�vʵܧl�;)Ԛ��ؾ[���ߦ�)�܎L�-�*�*P�ҩ�j�ʛ��Sv2��[�"�Χ'��k��)����|�ԃ��gu<�^���۷2�_�[�-�;��ѫ����d�U����)dD3�Vݦ�SM�d�]���`p����A�Hܔ݌BJ�Xm�n0?%�8�mE;Y�Ҡer;e*/{�;�.*w䡭��d�m����[鼩����ȸ�����{�H(7|�Z����
<�`��n�Y�K |󍤂������'�|�e�U��V�:7ڻ}��ڻ~:3͆���z��F8H�϶��Z��V�]������<=t_�]55o�4ɓ/a�k����[�V1�y��lBN��vj�ɫ�7~!���\<�J���h���������ɓQ�v��L������vs�s����ݫ���Te����9z+�]�[R�sZ���4���[����Q�8sZ]�e٦Kյ��'�W.ڗ���վ��|xh檗��/:�����t�h�a	"�c��Q�������C5U�8�weR�):��nj�(v��gi��Znb�[��BM
��a��Y_�*ȋ�p�k��o��E&#~7+r���c��
�~l�M4��ϲ�m"��V���%�[��V5���w�M�I/2�ʌ_�oU�~|m�ݗ��pߑ,��rI���G;����_�	k�E�lF~*&3-�j�H׵�S�Q]�N�i>�01:�6R(��g;?��hJ,j0X�ʪ��N���2��*�Kt�ls�t}�w�����נo�-7f���zuI��câ]yUI"���W����tFI���h��6YIc"���UG5Z9���}��sU^^�F����|����y�/<�q�R}��
���tK�/Z�2dɓ_vi�fюw��;�o��X����ͣ�v�4Ev���u��K՗�qIqIw�6�z)z+�;�ի��xUn�/.�4�<+�M���<)����j_<��n1��/���y�n `�*�_I��U���-@��	��>~~�����FzLr�N�*���;��o���v���j^�<5`q��v���F��:%�旸뛭�=�c�/kY|7j��F�������Q���7qڣ�F��?�sч��/�?���	�5|����S���?[�ӱzh�bJ�S���E?����S~ȸi2(�&:Մ���gۃ�eנi��RjM�x-�2(�;W�)V�ݶ�%��N��|H[e�i-�]�C%��Ϭc���_���a��ۭ�#�\�^J��CyZ��T_MZ��Vx�/�cin�j-���+������e����W��s�B�W��ȏ��=�G�+�j3�q�_D*P�Y��ZQF#�-�>V�%�Y� �r���VWE;-Y��)��H�򲛱|�k�ۨu�d���~�@�kiҖ�w�;e�������KQar�����Kf+���+{-�n�_�P.1�ȓk���%
ާ�m�W�S�2"|2�����Ir�ᒫ5/��G��ڟ*F�~ev�ݦ�����m؏�*U�N���26�2��&6
�����u�	ם�<4�Yc�G�N�`tKớF\���//��\th�G5[��ߎ���y�E�7�B@�������r�3����y���4��w᪚��ݚdɗ������
K=�}���������+�8��ɤ�<�^M��m{���E,�ϕu�GTɮѾ��L�������V�]� Q��L�2��/_V�[R����m�}��gm��?�A&L�zj��>�Q͍zr�jڗ���8jյ/w�D������L��p�H�u.VVm�}�W���㞊��k�l�%�R|0���q���8V����q�ʣr"�\X����̪�	�D�&����IQ��\�E7K/��Ih�ޮ�V�����k�r���H��,4m�I��@�ӻ)"R�eb�����e�d7�%-��58�ݘ=u�t�����id�t>�ݓFܰ(�6t���V{o�[lg��K�kW����46U�!rgӮ^r#\�sB�ng[�W�s���c���Ɲ&���ᓥ����	.����=d񖠺�E\������Ώ���)T��YI<7�j�L�6�	u�2O��G�r�T��OWD��uWD��V����yU:��]�}Wo���7��������D�|��T��:�ӽF�۴o�V�R�mKݣ|���Q�v����mĽ�R��.�WFh�d�O�*��I��BAH��d�{�y�//&�j^��z8j΍�]�}Yz)�c5}�&���=��ջaI������VԺif�M�$��w᫇�k��^^��F澗'h�E����>u�!-FBO�;�����2o��Wqў�T�Q]��/}�7y���Fy���ǚ^_5Y|�e�U�/~;Tsc��\v���V㝯0:?��4�\П�:�c��'��X�΍�݂���rP?-��~B�H8�F�'Q�om��+�,�Z�����"ܭ���ӥ\2�G䕑ۈ�ߒ��E��o㰅:�K��).X��/'%d�{خ+��T��샳��0�+�S����CsI�Y�	+-���q�T��ܶ�v���c]�u�^ܮOnB�Sr�͎&=����]ek����:�)
Or�ɸd�L_ʛ��[u�G/��j�n���v[u����+�e��s���n��PՆ�$�T�̊�ݔ�BD�~]����^��n��W��;i�X�����k}�ؾ�n��ȏ�y%	7�"M�)Z������$��C�݋�ɸ���с�RJ�u�-�޲?��I��z���n�6J�[(0��U@��j��5�<�����H���۲�wm���m����G;�=c"�}����]�=su��ca&�W��F��q�7;�z9����xp藵����u�WD�����j�r�㗗�͏��?7saQ�4���ǆ�{�����GT�e���i�L����nWɤ��؆��e�A��2��m:�j�Bmz���j�E˷~���¡�T6!&��@�y��_vs��5��������	�7>p�PR��ɯ&MV^�Ǟ���)d6��e,]oe׹n@�BQ�j�E&��`�I����&M}[�e��vwqѵ��Ŧ�L��ͥ�5�a3F�Ȭ5�j����B��`y��p�ED����n,�i����B��s�PV���ܦ������m7[���H�)W<
Jv��
�M����H[�m�셹INܖH;r�o%��}��?�vu�+]�_��c�&|O�-Ɂ�*�<����f/P���(K���6?����Yk�o�Ђ���F�����r@����� d�q��q{�K^6��aXғ[ul8pq�<�W���O�i�
^#���u�5s�OE��/*g�} HJ*L٥Q4�x9��3RBh���O&��ߧP,�Y�)7f��%���MtQ����Muq����J�%��ፖRu��^���U�޽`�muǆ��^k��e��vwe���V�9�\y�5����uvkɗ�f�6�}`n-c�F��y�u���q}٦MF��ޫ/GkWh߇;�9��'y5�n.%����I�p0?�����G߿k���F_k�jݗ�v��&���ջV��1ڻ5�'�},�=$m�y�s͛F<6��v��~��c,c~�Au����'��ty�vԺe�ϼ����B^����2&�獎]�^^�5xS.��'��訓&�뷮ޗ�:7Uh�՜������Ŭ�q�G6:��aњ_Fi~z0���	���'^z0�����>z0���������h�0Q<�#s��c*���dm�;v�N�7c��BY�c�ݖqH2�K&����*�i��R�}�R�Ҳ��G�ʩ����e7/�%Ie*?���6qX�ƻ�[�Yx~K/����;���d?�]�2�8'd��!k����T�M�K}��O>ʰܲ���2�J|��������K/
��i5�T�����v_�$��׭�aRVN۩�j�v[��o��H�9K�J��%��]�v�M� ����M�
��xk{/�.I6��������χ^/�ܶ�+z�V!��צ���J��+"���D2����ۭ�U�r4K>���!Y-.�K������k���?~���G��U�!b�4��K
�Hݔ�~Բ?�M�d�U�&)��8e-��-Y�I^�WnM�Û�e�Xz��A}��_����㤍����E�ٟ���\ё�|����Ŭ�q��q��8K�7��v�<7mK��k4�h���*�^M:7ݗ�:7΍�p՗�V���V��N��7��e���kkR�94^��`H�l))���@�G�!<��[���g���_K��o��o���Y_/�
dɓ&�9�  ��W0����Ý��m��u}}^z*ݾ�vk�&M/��5gF�8��vj�v;,��eٿr����"�Ȱ�I�d�ο�/f��GU�V�V�sN��R�.��a�����c|��c��F�9���訧FU�����@�|�_%c�Ԫ�JB��n`!- �W·{%*�oof<��YdN��+j�]�`�#R.�5��E�6ܛ���J���F�#��+n�.+��[�J���Xn92,)ݪ��TD�U���c�"�5���	�=�D7o)MP>�~�{*�����}�t��=xt���f������,�I��%�n�+�*>ρY�H�0n%�T�{p<����I��K'	����RBs��|&��N�U^dQ��7����/q.�:-p����T�����T���ծ��k�<���J��Ծ<+ɯ�v_��S&]��z+�L�2��&���y�&Mkw'y2k�oM;�hޘ�y�@�ã��Y����lmۋ����q��y�6m~愄���dɧzw�&My��y��]�Y_a'�����V���2e��?�A&�����Ղ����Ͽi#*ݸ����z�E���K�r��ʷgF�Ѿ����i{�W�F��{�Ug��v���V^���:���:�3K�s��Fz0�s��G�N��?�z����N�n1������z��Gbꍯ�|�(�/r�)W���X�`����,x����VW��~>//c��X�¤���cc"����b%��m�n�rˉ���;�~s���2��r��1M�S$o2Yz��+��!�cg�א�8r��_E}�R���B`V7-��io�kluku���f�o����򝴓vV�je��O�䒥m�>ʓ��a��#nP�k���� �e��/��H�X���%*��X��l��Ջ�P���lf|]�M�=���%o������9?:�؆�Q[�ֿ$�D_-���e�c�-�CaM�Te�}b��M�G�5�̮��퐷�^U2M�N�ȠY��;8q������~P��4؝�vϊ���r�}d��Kq�M*P��k���ې���˒B����;:̇��@����ϛ�ȘN���ɫ��D��Vr�5���XmQ����q�Dl�q�����H�6����W5�}y��B\By����޻4˳��N�Yz2�jݣ}�7���gF����2k��e��j_�d�ק/G4�f��U���<�7��������n�M��#�9�|�&L�2j7�vs 	�w�x�///j�\8a �����x��R�U}�';Xh���n�&M��e٦��󫷹���_�"�����Q����V���ExWgc��
��ʫ��Z�j��UR_^�����Z�4��t0Ѿ�2�j��Fk�U�X��*�<r(L9��xeU����:K%�|۸���ܲ,�q:�z���-��
;����K(�Ir�+Æ�~�bY��G���K<7ȭU�ǃ@ݰ�qSc�����r$��n,�N.�����־��&��[y��#q�Ұǃ;�������$9+�+v�K[��(dj��~hk�Vo��,<��4�pBD�2YU�;=	U�K�r3�������c����w3���)V�p���6ᄺ��ǚtm_GE�ޢ]%�r�T�Q]�v�k��҉vx�Z����:��S&L�4�&L����	欽ɨջ}٦M�ԺdӽF��5n�vi�aǙ}�w����G��ࠤ�ZU�BPϹ\����߆�����2��~�pգ��5h�G[�o�F��o�F��o�F��o�F񇞋Y�/�h��"p�Уw=zY���W�Y�I��2��ibdɭ\h���?�0U��l#Uo���=m\h^^�q��\ְѺ�u/u/u/uj���ߛ�2���v�:�mQ�����<7��F�:�������y�s��_�y�F62��'��H߸�Q���r�m\u��ݱ�׻�'W~�)r�m.�K^���r�'��{�^U>����)�fܡ����[u�ܵ?�%Y��8d�d�/����{+x�zv�"?�ᒤ���e)q�T�ɒ�J߈�ʃ�����\LD��Y@�a�M�R�-��M�ֶX��BP�RdP0x�u���#2*�I������)��4���,�}xn�3VB���$_���ǇY���Xp�y$�L�Y�S��c[J��d���"!����1�}d�%�[��Q�ƚF�צ��=��O����+J˱��e�*��m-ۘ�n䅗ے�?����K/�nP��H\:l���!��T�ƦF�JZ�en܏����{&׶��"[rL�n��[d�l+���#4�|�\�f���ڍ�c]��=�j�[��rt=6�+c��S�z����@�}Z�c>��W�I� n9ڵ��Y{�c��D'��`|�����BF�	q��<�th�Ϝ%ľ<8�����Ǟ��c����ݝ�g}��vto��F�Ѿw���;ӽ}��vwݜ�<6�c�/E5�n�D���W��RXɤ��1߆�l<�s�G\�;)
R��»s\hL�2ajՠ?��ϟ9ݻ	��\\'9ݻ��6�2頣#7��_��|[��P���8(���4�kKɔo�מ�}�+)o�aVz�<�����������5wu�]���vk�y�i``�is�����6��s1޵|������4L#�҉�/�'�Y�M��ҫ*�AK�`�9V]�L���R\X�x�5�"�u�GJO����בFK)#pl�������6P��N�&#�/!�d؎JJn��^U���-y"g�M��3������RYv��~�޻����	T��4g;v=sI���W�Rm���%S�Q��Xɶ����W]n���NA��c	���c�ТQa�/v�]/c/
�I�����yW�X�/"а����m��p��w�2Յ��v�3K�h�I���7���:3�(���I��dn}�����E�^uqݣ����Q(�Ir�.�����R��k�s]a_vxmK��kWݚd�ݚd�ݝ�S&���1��d�h�}٦L����/F�<8mK՗�V^�R��c��5\6�՗�q��Ley����&2���Wy���k�w��^����^���ݗ�v^��z7e��vwݝ�g}��vwݝ�f�:����	��z.!?��z^�d����662�&G�D�1�q��j�ExTo�q�G���᫣�;Z1�M�F8�v��Ѻ�u/u/u���Y��wE�=n1���q�6mhڻ:�U��/~luz�c������c��^��v���I�^�����'\������%���&���~�%l��،*���&�@��e\9X�W'�!|�!��xnvU
�r�U(��C��-�<���{zʩ�;y��.'��#H�6~s�.x�M�+�ҏ�e���+n�P�C�E����'l��Ir��2��&ܐ����+�ۈJ_�pUz����V��.�Ǜ()�&Kr?����",_v�%l ��e�d�o{o���,L{"���[����/��C��=��N���6��/���אua��Iѯ�AdV+�R�v�ɝ��9RDgn��iP�U?~J�����̵j/����졗��[
܃���p92[��J?����V2�D���B�o$-,Ϡe���f�^/���Ctߒ�Q-��ښ��K�[��ӵ�=�l�Z7J?���r]��f�~ˬ�g�F���@����n%��c���Y{�ڣq�4'�(��Q?�@����xp藣���tn�G5[Z1��ϯ�?��y�q�������;�����|��:7΍󼼝�ޝ��������v��z���v�����לǘ���}..Mz�Q�7���5s��olC�M'��2i��	�s�����F#-��Cc���T+�
�Si�, �r�SN��5n�y��������j]4��9򯱐WmK��ƛ]y���jt�Mg��/10Ql~E�*��4M$e�z7ջvԽ�j�/\F���ܖvJ���}�8-8Z*���H�0��6ܖ/��5uο���U�+^ǒU*������U׆U��cp�v2��kJ�����ˍ�,�헷g��ri:�q�g���0e�㲔{ټ�x�ۛ�T�!d����ؚ6x�(.�q��7ct*�
��*���2_�e�6�3P��t�y4b�T�h��/c�>�r��I4^ϯ$W3���sV+����U������ي�_2��z���r��W�Z��i@����E�=���.��(����w���
^'�(گ��>3�e}'nD�/�I��*��ï܊��(�dd���ޣE:��t����XK�:(��Ut�����Ϊ����/F_Z5n�M;�e�ѫv���F�6���՝��h�;ɓ_vwhޙ2d�ݝ�7��d��j�u�F��p�Ǐ��O���q�L�u2�������Ik6o0����Q�F��oQ�F��o^^^^��ޝ��H���,�`sy���|�0�����_��_VU���6%V�$�O	kF5٦��᪚�[��Z�j]2l6���F�ڴTn��Q��Ej��a�����z�����<:%��w:%���͎��;P=s@��q��luma�k޷�����y�}��q��E��Z��WG�=~L����v/��[���7l�����N��vS`��?�We;cv�o�/�@��rgn0i��n*nN�ʩ�d��Tܞ�.F䐫;��GnK)���-��'�q��(T����RnL\ND4�^�[8�f��s��'�j�J�1����̖�CM�ۈ��)P��vT��Z�R���ܪY��i����R��uҦ�ܲRxV�7�+���Y}�8�,�FB3�q;j2��^?��V~+|�MY�H[
����Pd�v�s��\9*��˨׭�i��C-O��I�������JR.�
���Ȼu��x�z߷;Y���r�m����%�����~�r�XT�#�>��+/��&��݂��4����^*�ZϒA�����b^V~�^��Iѵ�68N���<��Ǐ4�Tq�������H�߸tK��Ŭw��Z�qj_��%�\h�q	��$'�y�ǆ���������:7΍�|��;�˳]���o��g}�ѫv��v��ݾ��|�BD��Yi�]NvJ�i�4�0�̻4ɹ��I�R�.K�?�����4�����������^Mgg��޾|�I��\^/M��g��*�L�zdɰڗ����ך���+�S&U��F�<��~���!SeZ��|���ܰ���h��Ż*�ȵ���ޢ^Z�#w~�@���\I�sW����?6�*�^������[���ۊ���J��5�9�������Mݤ������p��r3iX��P�<Cs%�q<��VrU�U��k`֗�$�6�n�v����p6��vJ��O�����;��*Ȱ���,k�|V/�P5R����a���E�JLq�{��B�V2���g����s�9d�;�T�'>M�r&�"����̚�N��`v\M�b�$�Ӫp7V�s�_"ֿ���F�lu�lb$���F������$���X`h��KG��׌�ۓ�IT	JF�b�<�y4"_��Y%���L�yt�]%�z�����WW�7���󸂸���^uWWݝ�g}٦L���c���EYz7ݝYz8mKѫvw�z���L���4ɯ�4ɓ&M}�ݣ}4q�Ǜ6n}z���~tӗ�9z�<���qII	jըHHO���///////&L�2dɓc�q���=sc�u��h�磬dK��e�!j���ܷ$������A��5�z+�^��۴oM;�e�ѫu2j5n՗�;�h��_uF�9{�a���z����<���a��;�X�su��ͣ�;P=s����p=s\s��F���]�����6㝫��+�t�7o�j�h���7��w+=��~�M�m�q[v�+���m�ܱz�|���d�ݣa�	���ȐtYӤP��_;-�vv��]&�J/���QJvv�%wh8���^�܏�+zjg%;gX�bem?~˱�p�~��܂�o�����Yg�ɹ�@�������eP�.H�U^�����������2RE�gA�e����Ԛ����5��<���Cu��)K�)d�qyz�;
�֣nRTN�*���j~|gVǷrA��d�];i-�}ƶ[�Gix��)d��Z�?�T���ϋ�~��V��|rh�&##�Y*�@�����tY�,w��,��'�IYK�
U�%X��~ɻn��Q�-��e��2ڊ싒ˑ�XvS��~rS�;�ܴ����2^�u��ë��2m�~H���>�#`���F㝮w�:�����'��|��â^�<: su����ל%�o:1����6���<�����\�-c�/���N��N�ٮ�vk�^^]���f�|�;���tɗ�/y��?_K~!���ك��,����F��mK�M�
��%erTlC�"a///���(J�%���۳�tFRRb�T����H��sc���j��&L�<ѕ�62i?��,��Y��^K����6M_r�p��-�.+�jї�NxsZ����vʴ��Q�/=WT�m�u7JM�3��Wg�^�[Uy����e[ס$ԟ��;̪���"�J��g
�@ߚUI�}��V�>~T����tЭN-���(+n�U(\�u<5d,Z}��+m�86
��l#ڙ"� ���Oz	���0q���e�њ9%N���I��DJ&]Iqqɑ���sϯ�����s��VǝĚ&�YF
�D��״���M*�e#󔥎+HlcKBª&�g^x�i1��F�K*�mK��y\�l��:_�R�Y��_����oٳJ�L�R�=siB!EY=�2��q���j���ɓ]�Fv��]N����W�UR\���U�*����I���4sU�F��`F�V�BBBaÄ
4hݻv��v��j�L�4�]�}�g��j5n���X���j��cÇF�����V�sNy���II��8((/���W�>x��L�2dɓ&L�2k�����5sc]�F���H+�$�q�Z�"�ҁ����6�o%���wmK�MF��5nѾto���vk�ӽ}٦�^s��U�*5g�^�v���V��z���w�5qї�Wŭ9�h�q��\�`ty���5�;\�a��6:��F�㝬v�ѺL�2�Oq��_�N��K����E�-)f�7?�J���RiS��$X�[v?�Ȉgdݹign�Oé��b)7r�����[�ȹ56�"�!��l^R�qE���5kS��G�Y8�n~�.����;+~/2m�T��;�*B�Y�H\�{'j��v
�Vv��K4��iK�J�+�c]r,u���� �j1|�N�We�{����[ܐ}�,����E�1�Vv���r-��8V�����+zخZ����M�wy��{���u��C�G�y��쥗�H=ڌ�?��ה.T݄���ӹU�̔�����-Eχ+Zէ|���<����q'�uȭʫ�zoʷ����(n�3J��E@�kk�̟v���)0ƴW�+����I^�W��Y�"�y���ߐr8�~����ʐ�؝N�;[�l�u�<�}њ^ի�h��DO��H(��O�ts�kZ6��櫎��?:4�Όp9��Z�j^�kX���q�<�sZ����n���N��N��N��^^]���f�|�;��_Tɓ&M��#V�d٠n3@�/&^������V'}�o�O,��F�#))0%R����@���Ɗ���݁��_g"����J�k�,�h�Ύ�Uy㻛��o���{��mb����ɫח�@�I�$[��z�-ϱ15p�V�MF����
R��H����~:5`q��Fy���@ɣ%�nn�_V�_\utK��ǚ�z�]~�}�I�a�z%V(���n��Tc	k��I�a��e�3���g��H�ͣV�6/����Kʤk.�f�����e6; �Sk�՚�YU�R+��nD�ہkv�Bܕlm�ؖb'�J�a��qۂ��s4/������K���Ұ�쯾�C��{4cz�M����"�(K4i��&A���&iZI��nU����p��׸n\7��a���V����*�����,�Q��Á�Գ�;��9����䉰�ʬ-�8e\�N����%��f�z^���o���;S�ήo���Q.��&ϓH��Xz�]]�F�[��xs�4e�����//. ��}�իVw��ѫ/E2d�h�}��ǆw�&�j^�<7ݚk�z4g9��n�Ç�^�y>����zݻw��7��F�2dɓ&L�2dח�����e��f��Z����,��{"k�(��c"�&��B��۽�62)4%��	�_vs�y��ٮ�vk�N��N��^iyΪuTj�_�v���W�:3K��/��5f��U��j�lutf�њ_Fi}��c����v�?�h�/F��������5n���P0��l�~H��^!_���@��-��J��Y�!a����*����[���[,��S,��H�[+>ݖ|7{�m�y��ܫ��V��A�P$,���W�-�[��Cu���e���r!%BH� �aR.K+4�����S�
�j¹_p"����W$�֓���F���7V�ܧl��d��Y�A�쩛�VS�
���E+n˓�p�d_��)C�}:���b��9K�A��Ve�G{!����v}c{�[�J��9�Q�6��A�Gxվ�OVA�G�R���V9R�_-n�e8���q(w`�UNB�\�s���ň���nSv/E�S���JVZ��X�����k��[^*��òP����yQ؝*��I��u��!%kd[��*�"܆��c�����|��W��쳒�(z(�M�_˿`�4\aǚ^�8�ߴ�111��>y�ч�8�-f돟����	q��%���߆��<2�����VԽ�z3�|�N��N��N��N���ٮ�vj7������&���ѽ2d�mKݵ.�6y���W.���dɮ�Ѿ����kV��M9�KڵF^\Kڵq'/Vr�g/U2��ig�¿!)#W��o���6�l��lpdR�(D)��~N,~ng��k<�V��\֧v�sNwѣ;ɭh�)erR�"J��W��ի��[Xc|�p��W̽um@ڗ�E:7�я<�ͅT�D�n��5Ѹ����a�Ԃ���&ǻ^�@�ݯ�"��0�?�F�Ϥ��aGrO֝��;�I��іՔ���*P�Tu?*��'KFR���<k,���-�<��,�����?���Iڴ�a������3���Ǒa/�H�Z����ʷd/�<CU��<&�U���U�U�%N�r�U�R���p+V�6N�Ƚr�j�,�ZՄ��I,ߑj�x�$�.��cW>] Ȥ��.W;c$b�+RRΪ���J���X���;{z��:;���{Jm�;��j�Q;���mf��/����K�a�G�O���3BZ�qv_�ۊK8șgۈ�
��_�05UJ*��՗�v����v�۷n�ǎ�� v��ٴc����Ɗ5nѫv_Z��S&L�5�gV^��xh�?�=a<��u����O?`�$���ޫ/F�7�U-]��x�2dɯ/.�vk�U���f�5ٮ..(���ǏE��_>k��R,�T�/��}Y}�ή�ټ��Ȥ�a3@�K�ƙ6m�ջyj^��vk�KѻF��ޝ�٥旚�/;��F��6���WFi~z0�ц�:�j�w�z������W6:���͎�lusc��^z0��/ac����D�OI�®:��N�k���~�2hL��R�b�u�+/
��l5�a5�F��`B�[r%���M�P2��)/_���'��iJ��?�B��Ӳ���IV�w#�Mc�[�Ţs�o?�����^C����J����Mɦܦ�+�9\��ԕ���JF���M��y,�x,���;M�[��2]�+�-��2>F����)��S��X��L�IU��v;�I=�lE��V˴�|�[�Ʋ�� �7+{�L�Ƌ:$���죲��ك�X��d�N����gd��w�n���ۨ�ov�����;s��ʧ�����t�#A�6���+)���p驐ݕj۴�8d�FK/C��w�]�N�ʖ�%)��?�qS{���'e;�R���)�:_����q|p���|:B����[��)گ�����%�#�sZMk[���>�������X`ty�q����;����ћ΍��}�q�����^��jݵ/vԽ�jݗ�}[��&L�2dח�f�5٨�:7΍�M}�ѫvw�&L��5Wf�6'~!�%e��nV��U��2l9�_vi��ջF�ݻv�^}z���]�W�^���&U�j�d�?��J�k�X69:���*�5��6�|�Q��g,��5��-n
���<s���'��C�o�7>`Q�F����d�)d~�m�1W��%��Uc��.�qU��Ua�ũ|7z��XK+��%��&��'J����"�«I������/�b��Ȓ�\87��J��z��TU�l�2R��M��m���\�*�����Y�v�G�-�Y���)#Zҍ��!ZZ�A"��Gvv�o��\
w�&�;�?�@ճ��o���a��^^M�[���AK�uu���Ö����3�����`�q���ٕ��æ�v�2Шw*g��F4�D�s�[(o��yfT��B��+�I���j�ba��M�W;�e�kM�|���r�(~��{'I@�Zݱ�ۻ�:�\B����������Rs�s�q�DN<�q��иѢEa/'�Q4]�d�������������ݳ���&�Q(���-BX�Q�V�3��9�}�nݾ��9�s�۷�x7�N�+95�|o��<�1���:����k5f��'��+95��Y�r��۹j��I�R��e���j^w��Ѽ��tJ&j�sKռL�5���k�]���f�9ݚ��9�ƾ��|7���	��L$lg�Ț����q�=������a���D�֌t�1��4^U�}[�n�F���/���g;ӪK�/;��|���_�X���/k�v���/�Y|7j��/��un9ڸ�j㝫�v�9ڸ��qq�E�H.���k�[+_'�MI�r�`�l3��������ܿ���H;��&���ʭ���ە7[�!z4���(�*΁��VjZ�G�7=�ǢU
�JZڜ�ʐ��$�2xU�Ҫ<�Y��ߎY�Kw�R����I��'ׅIR*��[�����ܬ�M�Ǭ��)
��M��{1��YT+e
��rm�
A��+{"E��ն�R5K%�Rn�e���TC{���4����߶��$ݹi�vòP���n�;��/9�9�����)Ca �"���YO�ӵ��&W'���qeq6ݝ�YZ��ؤ��e�Y�Ւ�y5��O+Z�\��$_��!Vbڎ�"�'��pm�=Zn�J��۔��d�X�V��������e�~P��r��w*;@�VaY\N�Q�{iRnJw�ʬi��������~����m�O����ltRi[e.T�Wq9��VԾmn:��G;WsAD�����熎<4p�U��vxo����e�߆�[R�mKյ/VԽ5h᪙2dɓ&Myyvk�]���|��9ޫ/F��L��y|xW�*ݸ��g�*���y�����[���R�������R��^�/G�	�]���lj�S&��B��˷��Q���g}��#����r%���<kUX��w5ॖc`�7�Q���O8Y��`Nxq�Mv^�$B���ׅV"��;w��-4U\c��|谮滛Ό:%תڗ�����Ҍ��k��5�<$o$��v�'$�K;��V��s�0wv�����Oe���{�M62�����"�V�tܗb�;۽eY�E?i�J"?�I۞�󑝦��P�V�߳k����a!]��|�L�����u&k
��F}%���Y��]��;��uY�=c�_�������L*�"��+JO����oȲ��\���<m��6��,�K{��z���c�O�W��8�����S�	��щ䌧�,{���m��?_�����a�ȡ-�k�\Ү���O!\��X]�f�a��$�K��_�7��}l�ѯ�Rf�/�
�K�Ls����a������c�`�v2M/��E��jIU~G~�&�5jիV�\8pݻt	�s�� ��/@�緿��6��:��ҳ�/~=z������'^�sc�/V^�5n��_'�����q�����|5S&Myyyyy}���dɓNs_~<x�Ѣ���v����L��w�g�	g��N�l_W]|��y/w�O��5���j*)~�WR�������nݼ�;�;�h�|��K�j��]����+V����߷���_�ێ|���_z^]�52�ᗿ;�z��	���?sh�4�$g��	<�m]���RK,�\u'���_*ݳ�����BX�~Sw��U��J�gɦ��!җv�,䒤�9X��;��⸘����q���%j-�]��V���p��7g�N����:D���I'ܿ��L���M(�*P�j���l�;r����Ր��v��Cd�����[���^���_SL��^��cccr��I��<Y_���Q�%S5���o�'�l�{u:U��䡔ۦ�.V]F�/"��dT��Cc-飼lFR��\�{
���dk����E��\��s�jc���ng����6U>L���%GnZ��";��Em���m�U�+Ql���X?�R����.��M�ӵ�F���e���o*��qYv�\�SL��"�ʻqx`�d���)7$L�n7]��^�M&���_�g���Y�l�#�Yx+������?�s�//j�6����ͮ�q�U��z��՝�7|���qj�:��-fю��&��ޜ�9�s��9�s��&L�w�zw��9ޝ�ޝ�ޝ��^MGZ8j�ю&�26�dm�&WS��r�;-�Ν!H=~�M/��Ug_aI&�Z�q�2&��%�v��]�/V_��^�e��O�K9^P��������j�@��_�e�q�W�nJ�k"�Y�dJd�7R�S&�z9����`��ܿ;e[��P��(�m�L������1z�We��U�~�<��p�z��h����q�÷(lrռ�K�qU_װ��s�6]LH���R�K�;�$H��/����j�$+�Me�}�B������X��n1,���a~
���4e���܈Ī&
��'�P-D3Ҩ*���h��yC�����=ydC�"�繑�J�<e�l�<�j�&���ae۵�&�m���B������e	>����������V��Jd������]�x��Xn������f�Рu�Tkz��K,p�rl2���l���+�����¬dU�?��f�ʱq�H� ��ς�Ռ�u��F��_J&��nL�2��cK��a	I*���ȕm�}�F3_F5�K�*���O�O���j�Çl٥�����9�s� ɗ��__,�Î��U������r���Yk5��X�K��j^�[���պ�2dɓ&L�2i�L�2d�9��ѫ���jά�w�Ձ���a&��ϕqo��仇��}�h��W�<~t}������c����r�t��qk4h��/k6w�zb�����6�a*�uV�ڵ~3�j�*��kϜ�4UÆz4U���"�X�����Î^��n��F�������q�_Z�m1��&���I��W��0c$�s@�0sӗ���
�"�n
����7X˔n}�>^'��Sg���ً��l���Eo�(d��u�_i�΁g���d��Y>�C�����be���	B�<̻�`@���V9[u���_Y��J�n�v�J��҅gw!�,��F䡃�%Ct�Jv�[�WR�+g�XqJ��c!��r�(VwV����-�ʧ� �i?1��>!�׋�pa��47c���Sk0���!{x����Ca
�S!Yjf�//۩����n�+�(Vp![)g��!���2s����^��ǩ"��o�a��Y}�U���_YN���l��8��셥
��%,�K{J��i�}5f/��nS�ܵ>V�a�)D$�FW�!�8���ؾF܃����B��z��P87��(�ZB�S8�ڝ�i
�{qȷ,w(���K���<�mQ�Uv��ɗWmK�k���^�ڵj���/~{��N���`ty��F;�o��ޝ��s��2dɧzw�z����ޝ�ޝ�ޝ��M:7����n<����֌z:����� �X��w���/q��r�y���ϚHߵ�m,�K��YȳB������2i�/��F���Yȸc�|^wMe�eb�Ys��}�������g���m�ɴ��$���^&Y'��2dʴ~��rCh1���om�?����Q�<v���\}y��Ƽ�<}y���^�4��l����fa�k�ZL	4L���]l�dQ}�p������+� ��>l���ݍ��J�j$Z�WMM��h׳AZ���D�]��ŭ�>n*�}�6�_by0?�K?�ȣb��i�AḠj��K�X\p��ݯ�ߕiHP�H�=|���&�O��=+8,
�Ȕ%�ȡ��c��{)?�3�{r �[��[�u&<��gȭ�)�u7(mwY���%\��q~�{��<�v&���]nF߻i�������j�%N��ܚOY�qd�ryC�l�����=�(�{��<2k��*��_jʼ�ߑc�Zߓ}��FSx����
m���L:>����
��ƒ��4&����wE06��\@�����k�:9�ݗ�V�\x����<w�x��9�s� ɯ��/���n���vw�[{���8��L6��L�2i޻F���2dɓ&L�2dɓ&M;Ӽ��j����Ȭ��}�����H��>Eˇ?~"��Z�]Q¾�h���V1��x��d�7�޴yջ��\�^^�����N��j�F���s�F�6���w5۶��j�㻣E\٨ڵ}�W��v
��n�h�W����?>E���x�Z���8(L��1�yÏ�\:*��n9�W��u�W/�nF�*2E&���%�8��$Үؙ=��/*�խ��5�;��N�Kvˉ���P[���0���ݟ[���\I�%�u�ɷ��9/�,��B��W��>�cg�N�_�}Ī�V����d��#�A�[u5����v����������B�{XW+n�݅IY=Zv�U@�Bg�`l����>L^����R�$�E*P���YKd�ݷY��1	KM���k\knv�r�q4�W;Z�gm��U���C�
�ݻ���9V��FS��&��y3��ei�(H�q��!���R���=7R��T�2��=��ɩ�~r�:v�+ە����Q	Ca��C������I[�|���Y��T~�I�%-��sϠm0h/��]�/w�����82&�CV)S�����IJ�io�坕���n�+c�X׭�k�k|�]e�A����c0;1�����e��_uv��y�L�v�8q�ǚ�lusc��^��՞�v�:�ǚ^��5n���Ns  �2dӽ;ӽ}����N��N��N��&�V���֪ڗL�9}�`�5x�bؽ˷W�w������66E&����4�f~Dl�M�
��j�j�m�qnFI��>�h�	��'8/�Rz�.�v.B��Y)K;��ou�����o�"�z���}�6��`j�H9)K%���鵺ܡ��V-�zY�li �,c$���Q
ŷ�!
�����w��d��;Wq���V�\֮ڗL��kXz軛��z������̗��Uj���+������څJ�+�A��S��ķ*��1��,����ܿ�47VY���Yy<�{<�3�#���kn7�3�"^U	Ã������f�Z�_�c��'��^�u��r���&���o���u�ϗ���ő�VYד��E�nE|�����>�3Yő���� s����U�C#����n��enV��e7?Gm��,7(���nQ�K̦VY�����I��v�aK-7��V���&�$>����g�_���a��ʩ+���R{IT>�e�V)pȵ��-������YZd_Vv��V�^��y~�q�цҩu~:7tQ����n�wE����Uvwnݵj�>|���9�	�s��9� MV^�5gk]�_u;��K�MF��ڣ/���$ɯ�4ɓ&L�2dɓ&L�2dӽv��h�;�Y�a��ue���I'�dk�kܶ��;p8����\�i$���iVD�(��	4�O�"�Yɩ$�?�|��V���U.���^Mϟ<x�͏G<z1��V^�Yz5qѫ��k��Z�~l�sf�j��p�ի��Ϝ�����008�)!,��$�jK��P2x��jO�zO�1�b~脄��G�([��BD�rP)҆�[�dqG��F�Y���®�3FI�;9)�-�t���-����c�?"��s����7=)JM�g����/�A\�s�!Yh,�_�~ܳ�A��Y|��DL�?�N���ȬB�����/Ɏ�^?��S}�{�VE���B�V�)=�+"���nd�)ފw*;�N���[j�\����V&/�BߐvRk�o�~�^�"����{l��f&+�m���X��T����r�(V�����P66�R۬�?5���>E��S��,EjUX�Y�7�<�j�͖o�*��3�)Y!�5��T��[�%F���*���91��ܫ{�K8n�+-�ۈ�ϬA`� �b��g*��l"�ݝv��Y}�[�BJ���q��ɴ��
n�A�����["^/���@ݦ�r��޳'���9)�����0�sZ��z��h�����^L�}5sh��7�<��XX����V^��W�&���o�;��s��0 L�2iޝ�޾��zw�zw�zw�zw��9|5gF�Ѿ֌umK�]����������וk�o�?$,FJJ�gun\Vz��
�:�(b������_>�ŷ@�P)����e�S�(�+w��~/���-��Nؼ7K�rE���r�dJ���m�A��I�(��q�^mM��n��Ckt�6�����h���i��\���r���B�m��k}�xl�"U���v���M9z5sZ����z<����r�{�����X���q���^���r�k�e��Z?�r�xz�XK�ƭ���U�Ɲ����5�X�L�B��ʔ0�J�2T-��U������ۃr�H2�_�dCJ�O<�rz�{��3rH�p6�ll켒��$O����Բ
t�hɩ u�0�W�|�W��+o�od_w�nE�Ϸ�ˌ�;W5ă��/'qy�N���ұ�����e%7_�*M/����`R�=�<�m��~��ߏi�����u�{���8�T����gZ�4V$JB�
��U��	@���H����۱��_v&���0�.�n��?�E�_��&���$�%[���˳Q&^L�U�9z"s�4mZ�//. �����s��9�&L��{��6R�h�}٦L����V�Yz4j�L�2k������ɓ&L�2dɯ�;�o��f�ݻV�\y��h�k�5�+=-�*��ZL�-Q�2lHl7?ws�m$e}����O"�W��>�Afхy5WW��-N^����������FF```}����kXmK��F���*�諣E\٨��:�Xp�F��08�h�		�&&��zځ�����H��=l�?���Ȭ`�b|���D������D��f�o$6R��w!X��H>�fo�w84sD�08��,N�6J���\���6S������I�
nX��;u6��vUN�nb�1;�/:RCM$iCv2�W+v���1;�'r���v�9ȭ��$8V����n�;�`�!%U�^O^?���%)�J�y�Syȭ�����S�e�S��ܡ�²R6EY�@�`��Rn)M�M��ݣ� �f�ō�n/�7>��I_+d����H^�n�����1{
�g!���쥉��ww$��c�l�z ��RJ��l8v?�2��Y�;��2+m�U6�ʑV5�)�[���%��o[r���nܵ�N�Gd��v�%Vp�kϞ���䵶�K:E��7c){m�p�f�/�e���X���v�e�FJ�V�.���m�4�+��;����#�o�jdm�v籎��/G�����0x�n!4\\s�чڵW�]����yΪto�/Gk^`tRD����&�X�}��j��$ɓ_vtjݻF������� L�2iޝ�޾��zw�zw�zw�zw�U��}�ݣ~>y�活;�����`H��,,�-�ȅ�/e�J�\�
���u�v�_�p��9����Uٯ�r����ۅ~Se)C-��m=�G+YN��Z�[�Y�<��ѿ�k���ig��r$lbe��*ѓ�Y��t�b����]�<\;�����m˷�N�G鵺ŖA���ܐ��D���*�Uh�έ�|}y��				q������7sa^^Q.���}�wl��y��`��3�$�Hݔ^�-��6=���>���_[�QՖf�Ȍ���콲����FFC{�ʮ��ѻ_q�,Y��ߑI�)}x���IT��P��W��դ�s�v����f5��U��L��)���݌�@�����KC?�[�������(+nDl�MM�͟VE��RfÁ����?srH��-Ϸ���ѿ�g��-���"Y�g�p�.5=��؆?��^�DLd7_B۳���+]aRhd��'�D$�(�W�^*\������yں�2��o^^Q�V���՗я^v�4Qǆ��g9�ﾍ7�x�}��}��}��9�s��M}٦�F���5�gV^��7�L�2iޝ�ɓ&L�2dɓ&L�2i޾��5ٮ�9���ڵ�6�6�O���w��y�P��h�V�	dm���Y&��6z?��aaa�
�ĽY��j5f�W�<}yڸ����(�Ș���(/�=shǆ�{W�ھ��u��|��f������݁���
�dg�(.�|恁���9{UQ�6���FBW�����4��v�hН�,��>șf���DBY����N{m���򱈱�n��,��q]�cg�X�d�rD���~7%
gd�n��PvJ�e��!�*��;��ʭ��8�ҍ�*�R�E����O�M�ْ�v�b�~�J�ۈ��Sv���
����F܃��ed��wʝ��I_(�*F��G����Ws�����!oh;8�1M��hZecYOۦ�k��.v괘�{1�k�	��\��_*�~���۵�4>P���+9W#���)����re�X�VR��(u�{����{�C�Qղ�5l�IUoQr�Fri��O�zle�P�ܐ�.R�\��f졁�vV���ٱ�|G�0[�a5������Y�.,���l�#\�,��eOݐw���T&|+�˰����O�3�����Xm���O�[�,ߗ�ݱ�H;�ݤf|^���vy���V��|�0�������;�<�ڵ�\te��͎�8�.v�|�͏4�Tq�ǚ^�Y�M/��Yz4jݻF��s�	�&M;ӽ;�ݜ�N��N��N��N�i�L�_���N�闱��'���Նӭ���J� ���7��o�!
���չqm¿5n\R��~�_~��dn�p�h����_n�,�`�ig���z��ޙv������J���U��|�&��ҠV-�z�:��E�4��U���z!#c)%�x�10]~�K�̾j7h�v^����ի��h�(O����2.|��Yڪ�Et��/͆j��t�bw���AKɹ������v|$CV&�*�c�w>7�������_>O�e�����0�((Wb7�`�{��a�I��E�Mہ�$٠�X� �7e�ܴ��JX���Ҿ3��5��Y<IȠ���l���?*�ۖ"��l���������τѫ�����N��vpP9�2�o��Gr���*�`,09\���6�����n:v_����}$+W�����+
80)6k� �a��2�&��׷��s^?�j
Ҋ�<)�_F��h��WY�Kڵ�;�H(/0��q�hѾ��9�}�8p�}��}��}��s��lن8hѣ9�^^\_}�	�w�x2dɓ&L�2dɓ&L�to]��d���۩�N���m�:�H��;7c$�h��f�����;�z<��������y�מ�y��F�V^�����D�X�F�aǎ�l�z�Ç'���f���������=mf���*��/�E]*�\a��DLL$'8(.�~�@�ぁ�����mf��i<�Ay�����Xn�Æ�m��s�;s����5a$�)>��&U����s�pw���/�vvM����	�Y���k:�e�?��������S+��;r��nʻr��4e*�����TȆv;�M�]��D���e{$D���ge���G�pU*Vj�:���&�.E۬ܧ|������b�1�+)�!j)�h�ʈi���G��T����N�����շe]�v5�#�՚��W)�)F�b��M���m\Y�I�3�Y\�+v��ې�l���1Hc���lui����[���DR���m�iZX���J�qb�hWʝ�D6��.&�)Vv�d�m��e�z���Y�2�U��-L��e�5�.���%S!��T;O���A`��e��`�n�g���K7�K�[Rx�nW'���p(�}4�ʬ�JL^γ%z$�v��[�rS�:��J�n˫@�K6�L�m���d�l��n�F��Ci,�j��:6�ߣ�j���V�}��8�c��Ǣ�nr�����/����9�Q�.��y����kZ5gF��cÆԼ��e�ݣ}�g;ɓ&L�w�zw��9ޝ�ޝ�ޝ�ޝ��ݚd�mK՗��55jڗ�ן_�00P�y�n���r��Eᵋ,�����t�ȼ6
ƒ&��|���_g"���Q�i5�e��/�0(�ˋ�j���)ΝM��2�II����l�BAAX��Ȱ0;7798xd�vv�f�� ���j��їǆ�Ѿ��o�V�|<�s�_cW5���@��^x�i"y�y�ȓ�ғʫ{�_FvU��&�� �n�"
]�|�n���H˗g<�����ԗ-4�[��{1�;���'�yI��ђ�d�n;#?�IҨG�����IB���F3rT�֍'�x*N�K�ڪ�ڻ�Ci[��'dF"sZ�yB"x����tk��	u�h��#9��z�qV�7�1c�u	4ibH��d������oɳ�-��޼$6U�!rH��d��l4h��̓��>i�3O�O�	4բ�.��+8JK���K���h���.իk6iݺ\8e�ZիThѾ���.ݻ�F��n�}��}��9�s��1V�Q9�s��V���F��n�۷jի}�ѫv_Z��o�4ɓ&L�2dɓ_V��ޙ2dӻv�4v�;e�8��������ȼo��j���KK?����\B}]����*�J��! n..1ڸ�kF{Tnڣv�<7ma������}��HJ����7y�њ_���g��n q�@�U�޽my�Ϝ�|愄���ļ�Ϝ�10?��Ѣ��``q��������>��q��<8q�q���WW~?&�c����v�vy�V;۾d�#208��w�a��@����dP,��(K:����M� ��H��ݶD2Ԭ�owv˰Ҷ�y%N/�A�b)��n�nP���H7��HVl.}6�ً��D>R���E��d��Em�g���Cd��w�l��x��{Aۧkw��E;��W\R��^��Ȑ��F۩���u�Sk!z#սm���n�Z�d+��[�G�R;g]��m��k>۴ݐw��+%����3x����n���nm�Y8�v����|C[Q��k{r��Ca��B�ZVZ~����nq�N7�-cɈ�HY}��,��dCu5���M���"���v)BF�P6�v��m�*��D3��(n#Q�d�u��v�E�:��mMY�V62ʙ
��<4�O�W&m6�~�,݋�m�l�콐��7Y��IZ��+Q�M��$�F&K����vH6\�_?r�c&�͢��\>���63��?�y�k���8�.0��~kL2���Z�F�Ut��jά����ǚ�<ְڗ��V�[�h�;Ӽ�2dӽ;ӽ}����N��N��N��_vr�jݣ}�g�5�|5S&L�;Z1�ю�xHؙ4��Y_������2��
���7Ksu2eZ)�.ޙ2���bbe�)x�cc{aP�˕��o���6{;���D (����о�4�.իv�P����n<�����2��}y����Ƅ�3�	����^��n|���6�������a���4�(�$+�6�ry��M��r^\f_5��n�cѳ���}�܂�qK��.6����3j�U�B^����&��bȁ��q�cj�E�n�:I�u�וZ��ѱ��Ep���FYy8vX��֭"&��mF\������sK����ʤ��*J��QZ�/{�<�1�{,`v�n(�*�4B�6"�g��~l8+�<R�̔^3�=a���l'�8��*�k�9ʢP�p���i̴�i/��ҭU�7�}���V��V�Z�jթ�s��9�s��9�s��;����9�s���v��4h�s��9�s��9�s��9�&L�2d��|��|��|��|�4ӽ}��vwݝ�g;ɓ&L�2dɓa�j��(L�7�1�͎_Fi4�?w��Y&���~�曕��Yd.���{|T
6A�l��﵇��6x81���1�}�ts�v�Z6���XXF���cci%�n�!#c%Y�񴑐���Fi|2���<x���/qq�����ի�f�Ϝ�^������o>sKˮ.0����[Z4U���		�&&�������;�y���4ܬ�+� 鵲n�n:M|�C�˭�ն�W�϶��X����!l��jn������em&�ŋ���BiH6����JU�F�JR�W+��ݠb$hT��䐽��,N�/ag
�I�r�0ݝ�&["����l$��fJ�"�����Vݍ*���/��e.z�Oo����y-��v!��*r?����U3r����w��� �,7$���������}������vU<�n'�B��l�u6�J�����2)�}zn^��5dk�d����"��ϊRݶ�u�/�dvR���)#���W9�~}b��������ܱ�asݲ�uk~����&D7S� �j��w%.���L�����e;$/������d�[
�K��qH;��f�=�vBȈg~��+��[r&��L�C�,�e� �pw�	Kg!�J}���r����i��Mk�!��k�wxe(<1�b�-a{��Q��[��Q:?�Z�qGi��i�3��ڵ^��.0�˥��|����Y��w6:�3K��/F��^Q�u2k�o�V�d�mK��F���hջ}٦M;חf���;�������ӣ}5h�v^�5e�ᵣ�˓������ɬ�����
s� Kڴ���II@���\��y4�E����ُF�{V�{;1��~�X�����hNs��9�s��9�s��9�s��9�s��9�s��9�V�'�(ؙe�����p��	kF?�I�o�U�1�R-)R^��U��a:���G�!k2��?��j�IVZv��ɋ�d\[���Ǣ��M�=~��JA�X�9*�K'gݣ�cݳ��9�Ü'ez&���X<�b����g��L�*�B�'�Z������hKJ��7X�n��'�n)3.':L��Q2����q�&�fX`�������^Q��ta���ґD�Ȯ2#1ʿ�G��2����^�B5g.��cj�rOv&�2�NgZ.�_躺ȡ<�A3�`����j������:գU}�3���V^�۷g9�}�hї����������9�s��9�s��9�s  /���s��9�s��9�s��9̙2dɓ&L�2dɓ&N��g}��vwݜ�&L�2dɓ&��5��u�	�&�O�}n(���62���Lfw~�H�3�uu�$�hl� ʷ7%���y�P���ѣ9��۴o��5�Z1���D'�R�y�����D�W��	���*��ͣlumZ��T��ի�f��5x���w6j:4U��^����|��h�׭�>ss�/��Z���<wo�����n�cѣ�[]~�ʷc��L���c��K�~J�W/V�r��U7+���rҮ(��/%S���iZ��i�=���q�7n"�@��x���v�O����C%����U��g�%P%,��;c���w%���6\�)��� �e*��۽�D6���RJ�[.X�l���)�}����I*��n�t��r��H�bj0�^�V���7ky+',ݔ��e,�Lgd�"�l�2��ܖSvR�!��f�C���|��[�vv;+)�*��+�qIU�.§�@�NU��*����BnQ�«�I<7ggm���iZT�>�Y��)|X�~��I�_�o��n{����!,�JZ�}e�A�HZ�|+L�D9\�VSo+L�m$:w�+�rA��b�?rW��w�~IK����2v;����;� �k��֠pp��Q����G����8�5ʷ���Mwy�ɒ��dl�o+�;�N���5>d�)5M�[�a����$��sBZ�q	��߷�����=`j��v�6KX��O�:<�(����08����D�Y�5�_5Z+R�q��V��F��ɯ�;�oL����h�V^��o�4ɧz���ݝ�g}��vs��4��v^��z7ջv^�[R�sZ�Ϝm���U'�I����F�2�����_ww�!��ቍ�E����E��܃ ��
23<����ߐd)
� �6x8"s��9�s��9�s��9�s��9�s��9�s��9�2d�պ�4$O�O*7��я^k���\�\5�\�	ab�5�F�3R`I�Qx�hؕ���t+��ev;l�%e�}�e��!k6\��mJ�iE���%�-4��(S�a[������Q�����3 n��e�,�|�(���:2x(MyWJ��E_V͇f|���E��Fc��y����N�J(J(K��(�n����,�ߐa���+��뤽��άd&�dg9d��2E���%E�z�B1\>ʡ7)ܟeT��U��d<84��Æ'f�|n����Ҍ[��^��z4U�j��/N�Wpڗ�F���}�ݻv�4hѾ��9�s��9�s��9�s�� 9�s��9�s��9�s��9�     4�_vwݝ�g}���k�������;�������5��7�By�������_��V010^bc#+��V6�t}����
O_���v���RK$����V��>a<���G�l�hї���ׯ>|�d���6�A�e��,E��Ύ;V�9�vtj��6�_��1Ϯ�~�%�㣛�4U��_�9~|��h��5V�Æ}zځ�ǣE\x��������H�th�}�8�Mq�E���r�~S�Y-��/)m?ɸ�4�	+��>��,ݶ�iҖ��?)@�g�ҁ�p�ȏ��b t��W,����쥺޶+
�S6�)WW�~��n��g�!K8��nw#�J�qH9�}�ϷM_�%o�R6�)��`ݕv!ʐ�T�>w'��d?�K�@�W�S�%�05�)ec�?������P�?d~'���l��ۆ�)�8nKQ��`P52�ƶ����j0ݝN!���64�R��|m�5v��re�[zj�YZ�2��93RrnG�����榿�;�[�2ԭ*n&����+��n�l핼�K'R���7�/��E���3n���[�սe?�B���Z��"ۭ��0���s�E��ͭ@�H{\�{9�Ǳ].�vB���K._����$hV/�_�N����m�fCo&/c�m��;,�+'C�"�s�����"F�D50�+'ۋ�c��}�B���,zvF�7�e\�o��/j֌���p��f�W���Z/���i�4�h���wy�Q͚��W��W�[Y�Q��dO�0:3c��^����юԽ�j�L�w�y2k�oMv��e�ѫv��L�w�.�F�Ѿto��;ɓ_vwջ}[��|��v^�[R��l�?���֌����_zs�۷Ѣ>�s�uaT
*�@�۹a碎;Z�[�\��M�1w.�>���]���=�w)C����t\\Ns��9�s��9�s��9�s��9�s��9�s��9�/�Ժly�a�kG^r�,�6�4�߇�kW&����b�l�M��n]�ͣ��ո��Ƒ�O��,e�"R���Fɰ7xa\��F��cM���r��Y>���rdV���ϷVB�p�e��˲xM���.�tg�}��W�v��xl�7�}���2ͽ����>E'���Ij�
Ee���ܗu����Q����{�4X.L�{-�r�בU�p�ko�5����3RB%˃�ܨ��c��/�cj&���Ԑ�Lț��.��ը�V�r������͎�mn��M�5�yy{�s���}��s��9�s��9�s��9�` �;�s��9�s��9�s��9�     4�_vwݝ�g}���k�o�F��o�F��o�F��o�F�8j��������1?p���2'?w�Y*����\�>�X�ij�ij��2%����V^�N�����r25�wp00$R)�>mZ��Ϛ�p�:8�K��a"��b�.>�??n�W5����֍th�qW�/��������j�4UѢ�>r�����W6j6�_j������6j4h�`q�������e��Ǐ�$e��s~?�����Ekn?���x�k=�,&m�cn��3Fȸ��W/�{����n�nJ��V5����Y�e����f�/Q�e�\���E�~�+��b������u�܅�3�8(̋l����^��-L��I����զ�rYzK�]�e�r͹
^'^��#�{��4}޲y���/	&��ՠH:�>DCWnB���eL�grp��'�M#v�r�h�O��rgw����v)�(S$�����oMZ뻋�V��VN)�(l$�y-���v����R}�6�Q@�[���C�v�s%e7������$�c;$C)BF�i��]mF���)���n�^۱۲��%OJ�� �a7l����v���ڟeoe_� 併8�[)*�r�Zgecg�X��J(n�����!`p����mX�Zۦ��Y��ݑ��|CSm�֣5�(�ʷʭY��V9��nƁ[��61ݸ���&z����ߏ4�c@����G;�sN�6KXֱ�:����Z��_z��``q�g�W�F@���F0:?����U��v��;ɓ&L����ѣV��f�4�^]���|��:7�w�&��ѽvk�ӣ}�z4e��\\u��<k� ��1;�q�ћ�:2����n��Ksv�X��ܸ���N^�n��F�Z��W6?10^b`��.��9�s��9�s��9�s��9�s��9�s��9�s�}٦��6>y���2
��e��эV�����~�����G�-��K�o'�㵆��O�����e���&U�ǎ�a,,%�sNi͏��`�p0!\6��<�x��+��J۱����g�	�^��'D$7V�+��&BZ�'��cj��r�X���cM�&O���'�����J�7yd�䪯d�F�؆D�B���$�p�W��)J;+�,�q�������ܖ\��0k�d��tI��و&�!Am8]J�.��*������Q-_<w���4l_�.�a�����Z�ED�V���~��q�V�֪�Ѿ��zw�y2iޝ�ޝ�ޝ�ޝ��s�����nѣFs��9�s��9�s��9�     4�_vwݝ�g}���k�o�F��o�F��o�F��o�F�|xh��j�Fh����gk�Ō�Mag"��;���&�҈V�u�BP��d+H�^������Z�PPY�f s���L%�M�}�����_���U���GGY|�$Y0Q?�uϜ�;�07a<ڂ��	��ū��q㻛5*��/qq���>r�����W�ۏ�n `q��qaa		��ֱյ�����Bu�/���>F�C��ߦɵbk�"pwᲖ�~ˬ�Y=��6�T�ʲ"�[)[��|�\��//
����حo[�����?��V���_F�o[� �s�*�&�Ƭi�0X12.��BY�!`�3��U?���}�8��;���6�,^�C���P��^ۖ�������'��g���~Y�@�܏�H���d��$Q�w(K��������)o�[����V��oZ�Ր�}��[�a��Um�����;gQ��h?�&v�*��t����*�m�Gv�(T���ݐ���f�Z����R>���J���[��+~ؤ+S!�;ؤ���v�C�ᐫ2Χ��E;��bC���>�)e������94BOr��q8T���G~>1O䕨�v�����Ir�(��J�Zjvw�e�n���ݔ���g�2�*n�^r7>���C���(�V�� ɸd�i�u����{��)�]EoY����2M��D�w1�F��K^��֮>we��]�U�\u���<�_V�/�tY�)$��|�Vr�Z-Q�l7o�_Y|5hջ;ɓ&L����ѣV��f�4�^]���|��:7�w�&������L�zto�ϟ�����;�s��0��}�ݻv��2d�`���$����L�G�6r*I4�G�+��L��9�s��9�s��9�s��9�s��9�s��9�i�&���xnѾ_�ִcL�,����ȵq�Fx~�g�\�eR�p�<�a ����)V��=�N��'��Y~lk��}��'�^Kѫ���^3�Iuc�����J[F�6?/c�Mc	�����HP�81(�^s���Rv��dW.%�K��q��lX�K�˹˺�K�{{;u2U��'�����*�_e�`��'�������`o���'��������Y�Z��j���dX�d�V4pq2�+�X��)u\�� ���TgvԽ��l"|�AQ�����]���Q�/F�Z�n��W6:���ջ;ɓN�dӽ;ӽ;ӽ;ӽ;��}��9�s��;ﾍ4hќ�9�s��9�s��9�s   ��9�s��9�s��9�sM;�ݝ�g}��vs����Ѿ��Ѿ��Ѿ��F�ɓ/f���������XX�}��������k�o�����J?!H\�T�_W#W>&2kQ112i4�667�^�q�Mv��_puu����>�/�̉f��^A��`��q��\tss�͢�y���4]���qV�5]���W�9{��008�����hp08�.0����%���l��}}|M�u�BXI��x2�}}��(U�$f�~6Mr�&�	"��H���~��#�d�d&:M���+"/�խ�2�6N����DVB�P䬼R˽���4�n�[�z*p����tވ��YZ�ې��R_+��J�x���e�²��n�[��(1�>!��6��J޶Or�щ�҆�bVÜ�~�v�q,�Z���g�a��I���r��vӢe��!3�l6�)8�u��>J�ǡ�J}���l�����/ �V�{r�N��kiPą�V=�L�#鸛��7i�[�[w�X�Z��V�������j?��g�Z�oj:�O#����z����eg�Z���C����ocC�e�R*�N��{��D����|ʢ�$ߝ��(ld=�ow�A��E�]�]ov��Tq]�k�?��Cr��*޶Yە�o�{-�Q�F�F�ȿ2Q�U?-��V2�FGn��m��8��ݠ�14�!��P2��FNR�۴��V/SY��s�|�����`j���G^|��n*��k��<�e�u����9�VҎ�Ƌ�㌂��9y��/I�Ya	q��Ug���ګ;��km�c�;ɧzw�&�F���hջ}٦M;חf�|��:7΍��ɧz��4ɓ.έZ��f͛54g9ݻv�7�|�9�`	�w�|��U��vxe�)#p5t�k�'�]2��͏�lf~��$Bag"K�L��9�s��9�s��9�s��9�s��9�s��9�r�j՗��6�y�cǚ���*8j����d�V1�:��V1��s:�щ��~��I<e����cpl�)��u�E,f���E�x�o����$O�4���	"�N�U
����*��:$��0�T�â�Yqg,�*���I���,xuQ�����&���F�<lٙ�K��w�}���W5�?�%�i7��cS����ͻb�������v3�߻I�r���M�կ��D��}�T�D�c�<7旜M��D���J�$�	��q漗�v�x�5[�f��2���tJ%�ݾ�ڲ�p�/F��L�4�&M;ӽ;ӽ;ӽ;ӽ9� '9�}�nݜ�9�s��9�s��9�sL�2dɓ&���;�������;����M;�ݝ�g}��vs�������;�������5�΍�sZ�ן��--���6�
���]��n9��$�\=���N��*6����ag"������Խ[��Z�/F��� �Q�Gj<�����\�Z]���C%������p��Z]���.�u"���qGf;L�����G��{�������HNp���!9���^������Ddg���M&�����8g��w$�y>����e�ӥ/�U7�r�'��c�_v^펕���^��	W}�M,�����2�|F�+�@���[l�Y,��w��۔=��4�M�����ݶl���VN��!{l5�9���r۬�e�8�_-����Y\Oe7[����Z����W?c#C���(,�l����b2�F^/���Su��?.����M�'&M�Igr����7>�'ݐ�c�Md������Z��Gm�(�}���[��gr��+���?4�F�VH��R�u�;<^_˰ϔ��m7g]�Ȭq[v>�~���D9Y���n�C�S�r�&�H{�N�o;������W;��j�2�E*!���b�r}�4���M����"�]���@�n~gj�dj��V�d���!��+r���)C���~jr�(nZ�J��[��忍�/v����6M�Q��ǵ:�wd_g��C��
��J��J\�^�7;�N�vӹQ2n�=��+Y��q2���k��q��m�󸣣�\�2����q��9|���|�����������Wp�c��}'��(�suц�4��i}�ᗿ�l}`n4s�}٦�F���2k�o�/F�[�ݚdӽyvj7΍�|��;�^&���Ѿ��L�2��4hѣ9�]�v�ۢ�۠ ڵy��_*������܌�K),�Vz����m,��-�����	�'9�s��9�s��9�s��9�s��9�s��9�s��N�k��2n��n��^^L���k�O9�n.�a�_�5�Q�#pl9������F�d+����vC#2$ݶ[l����\��j���~!�ɹ�OI@�$(V.�q_cq&������X���</?���R�[��ߎ�o�m-.����i)	�ٳZя�l%_6��4@Ƞ�����8�gı�����r0�ZJwO�^��5����к^]/AW�XI�j���#q�Z6���;�V5Z��3�ۺ1�Q4a��|�*��,���	/�Ddflٯ%���bbb`�aǎ�3��2iޝ�ӽ;ӽ;ӽ;ӽ;�  ��9�s��9�s��9�s��2dɓ&Mv��h�v��h�v��h�v��hޚw��;�������y5�g}��vwݝ�g}��vwݚn�i%��{	F��ܫ_V��&>�n9����dg�o���o�nqdvk�����O�JHț�&Ç
���		/q�G�]�;��gm~�X�S�4�G���W�/y�j�������������23�dg����n:��ϭ�����я޽m``W�i`W������0�W����+������d[��y<�v�J8bT����b>YJ��7S����[�)U�O��BJ��8�+��IJ�����l��j9l�.P�[#u�}e���>!���Q]NN=��%v[u��x����W�m�v��r����3��x����B�����)l*4Mg-$G���o2��$���W��,2"(�Z!|�8�������Z�n�;ɕ�ɣ��yC婥m~Q�Y�e������e����rW'��j1��RP��ڲ��&�z!�8�o�S�H�^�VϊR��i��mEÈ�D2��vR���_l��S�!bc72����ܡ#J���r�������Ej�vR��e�98��/S���~B��d��v+}��K�Y鵱�(�v��ñ^_�]�Y}_e#p�=����Ȃ>/����~b�19��W+"�a�P$���)�P2��}d���~IR}��%������o��Pܗ�M���ß�+�����;X�9��/���Lp?�y�端"���ם��������5]�ս/u����-Q�������k���w.ѽ5�nѽ2k�o�/F�[�ݚdӽyvj7΍�|��;�^N��7ѫv��&M}��s�V�Z�g9��` .ݻv���wnݗ�j�!Yb��ܫ�_�lgX/���s�����r���k{p��9��E��U͍9�s��9�s��9�s��9�s��9�s��9�s��Ѿ����Z�F���4&�q�2l�7���皎<,�]n�հ��ϓq`Q���5����+9|p_��u�&�ߦ��cn/�N�b�Z��X�ȳ�"�Յv���%����U�ھs�+�M�H�[�Z����`q��Wū�=s\h�њ&¿o����w�``p�V�?:%��K�)<��F0��n���B�)%/�V��,������_	;�+�R��^xפ�+	e��+ʯ8�n{�?�t������U�^����6��Z1�*�����O߱�UmK�MV^��z)�      &���L�5�pڗL�4�Q�v���o��o��Ӽ�2i|5SK᪙6�y��<6��V�YyypZǅ5�y�c��u5Y{�c��<��i?%ˋ��_,�cѢ�Z�ᗣ//_g"��EX�;�B��223kY�cMv��:��T����7���<��,?�,�.Y,�w>U��F;�X�K��W�[]zڸ���_�Ů�%�3U�^4l$gX(�`�BAu���^~tc���������G�\q0�����Ύnr�y�c��ZH(��dXpę�R�]z��>pY���nl�����&~�']��%���WiT++�%{wk{=�C�� �vr�^�%�ߚm*��%��V�u8������$���P��~R�1%|��x�T��)�X�e;����5�rh��SZ��+Z��$�����D��1�����u�k㎔=�F&��e7�n}-�)l$��V����^�w�M�V���ܮ%�Y�U��d�w)R��e���s��k4���J������~����
�7e-�2R6K[o�bb�����ND7�˭�b6��v�s�N�`�k$[�n+o���c�(`��p������]��n�����{!���w)@����K剧õv�|��*�K����S��,���$^
UĿF��Y%;��W�2��J^N���%I^�n>/�Y�!oe�{-��������o���ܤ�,�/iJ�64�.��F���͎����?q�Af����8(�q��;{z�)����X�����O'����͚�l�q�j���_��٨��G6j5j�ޫE�]����|��v��z����ѻvk�˳�����vs�9ݜ��wg;������vs�9ݜ��s��;������ޝ�ɧzw�zw�zw�zw���ɬ���i6x�s��j�>a!3s�;�@    Ns��9�s��9�s��9�Æ����V�۷nݫV�d�7���W_�vU��c*�<�y��O��w���rk汉\cf��"���׈~Z��N}i)0��_ٟ�����*���`�$�^�)�ݬCdܜ^p$˪���z�]�̽$m�/�r��/�y�f��L�i�գ/.�;��]�k��׼��`�dJ�sѸ�;r#k�nRz���o]��b�j����W�\A��DL���:Ie|$O�}y��Ǐ��$OX�*�t1��6�Z�l){��{������/��(L9�_V�֓_V�_�4p�L���gF���     ɧy2d�h�/���(Nw/�4ɓN��7ݣ|�&L�2dɼ�����_vi�y68hѣ}��}�&����h�j]2nw�y7���4}����W�X����}�aǎwn���ϭ�6]^���M&����Yd�O	�֌|�����1��d�燞8H�>F�����[�m�/a'���_�[\����W�[P08�����7���	��\~n-@�U��W�����`��y���
���oQ�V�7��ǅk5�_l�8�m����%$�_n�vQ2�;=�~�l��oJ�N�b,u���޸0�X�v:���Q���72!Y(n#QY�g9j�S�����e��.ܖ^�s�vq�=-��g�gc���dd��M�D�b���d��Yfܡ��o�����d�<Pܶ�B������l������S��Ir�;)��{o����+�N��r���e�F\�����G$���'w4��!���|����J�[u�E~ܡ'ᒳ�4:����k�^������̮�.��
����r![�JH�����ln�7�^/W�_����V���4�+n�/�����#"!��ܲ�Q���/'lc#�-�e��Yr���>J���U3n?��re\����a�&��_��Ҷ��\�(�s������UN�ou8�J��c�V'nJ�צ�2�:ճ�춭X��rnLܖ#QC�Y{���o*H��s��V���'�Yx˕��U�(\Ri'�V�X��8a<���/	���~wq������o��@�ぁ�����<wq�j��p�ڵ~<wq�/.��Q����]�/Vx�Q�E/Vxj��V�[�ݚ����vs�9ݜ��wg;������vs�9ݜ��wg;���������9ޝ��L�w�zw�zw�zw�x]�w �Nss�۷o��   '9�s��9�s��9�s��ի�<֭U�v��V��4hݻu2dɰ�Z�dH�U����J�wp���_v2�7V�7V�^'����ku���)\X���	F��wT[t�lC%M��ȓ\�5Y8�����*F�²X�*ݶ�}%��v�����h�~�Wsa����7�^��۲�c,c`�bn�Ѿ��|xgF�ʷj�Ǉ��ګ�
Oݤ�q7l]�a��ud�t�d�Niy��7�������������f������l�JU&��������/��8�K_��U]%���kkUmK���vi�&���<3�zeٮ�2��z      	�N�dɧz�[����>z՗��2i޾��N��gv��h�F��5n՗���Z5n��V��^p���jի�n�/���MV^�m�_V�οť��S&L�	ݻv�[Y�@��ǣ�m�����X{X�����D'�-\�e���LL%���Id�_W�����H�����%���U��f�"�����k5�|����F����٨��w6�yቄ�������: �3y�kϜ��u����<p9��Z��v��3K�a��E���-_�5~���M�irU���$$n��#�!�����,u�n[�-�D1��rh���4��ے�␰b��n��B�qH_.�/��P���n�H�I^�v'vˆ���o�Y=�^�Y���ܲ����n�Yr��P�7�����d~I\������E�;SZ��d�C+Y��V7n7�˹e�~b+4�*J�[5��7{���B���ݹJ�~J��S?��dTN_��m�ߒ�Q~W��-o[ײ�q{����G��:qM��o�m�nK��5=Z��vA��u4�nZ�*�j|�P8d��7c*䐥��}��K�?��퐰x�v,\�۴ݐ{��*��h*���"���[L�����;;����#�7d��0�]�Z���o��Y�����U��d���M��R�-�Թ$-��)��.+�s�ڏ�I�<Vxd[r��x���D7>���Y{��Mj������}��P-�h싇�Y
�B���6�O�a�q	��G>r�y���O2�`j��]@�㄄����*��F\x���vի��3�j�x���w��w;�h����ڣ	��^��޼���vԽZ�o��9ݜ��wg;������vs�9ݜ��wg;������vs���;��w�zw�&��ޝ�ޝ�ޝ��������Z�k6l�hѾ�����ݻv���`  s��9�s��9�s��9�Ns�v���իF�8j���VԺ���o:#d�8<��p)/�����^�O��m���[����rp���^���	ga��ٷM��[h����ۤ;�S[L��%)
R���YK>�������/v�kWmK�]���s�zj���rk=��n�vz9浏
d���������)fm�5^I5�)4�k�($e�;�"`tA���,������߉�����~�~�"�ϸ���&�������BW�a�p�{�˯&]�5n�їǆ��{���q�vk˳��&^Ú�     dӼ�2d�ݝ�7ݣ}Yz6��ǚլxnѽ5�gv��h�}�ѫv_Z5n�M�6�i�ś�g"��\u�'9�s�}Z�hջ;ɠ|��q��De�Le�OXK��((؛�O::�q��^���Kڴ�u}��1�|�&M;���_,�y�q�5���2��6�O,�Ϥ�J��P�V��&�^A�{dlF��(e�r�we@�Sn<���v�Q���F���_�E\x���/Ϝ��j�tK���	��_��As���Ϝ�����6?8�藣j��\��a���p<�h�/q��'�>~�ݶ���`k�e�ȫ�����Gnˈ�~V5:"t�.R�ܧlt��؞�^�d*������$��ϧl���?��+������5���C�[���L�_�%@�[d��lV����ڍ�[nA�b2��*ov�Y
�ݐ����BJ�v�[؄��ۭ�#�\��7����6�-X�ӒB��V��r��"�c�)I�4�U�n�/۷��ld=�)��J��j�}���)�N��ȭ�u��2�e�qJ=�Q*�|��R�݊Yq0z׻�(S7�Uky���)�+gJF��I��=({j1FNJ��켪d*˳�ې|���_G�����[��}XnʵIɒ���o���#�Mr�le���C-�ɕ�	�	c�a����	�n���w�f�,
��8�2��mw�9�#�ğ����a�eϠe����N�����7�����2D:>/��r��e�@��d-����TnU��l���Wk�F^�@�Vb�lLM�����_<<�h��>z'׭�`j�u��⍭�dI�, ��ͣE[��008�.0��wF���Qǎ�<wq㻏�٨��W�9{��<����v^��a��������yy/F�z�o������vs�9ݜ��wg;������vs�9ݜ��wg;���g}��vs�;Ӽ�4�N��N��N��N�4nݺ�����r��ۄ���ϝ4@��v�۷n�  Ns��9�s��9�s��9� ����ִc�ǅyyy{Dg]�q�u\U].�-u��Z�f���û@�Fʳ�\�2�Nt��;�S�ǆ&�B�rV�����5�&�v)l��-�P��4�<���n#$эz�5nڗ^L�v���M��G^i�z�<8mKյ/��d�۹������'�ݯ��vX4�R/(��w���h��W�����H܎-˔+��E	c�������5���X�``qvAH��࿭UZ�&������;�=z�������`}�����ɓN��e�&^��     i޾��4ɓN�d�ݞ<֮:�ͣ�7��V�Yz7ݚd�hޙ5�^z��Y��hջ��7�|��BB\\\K��իV��Zя5Ɗ�4�M�"��2�7^幹�����g��������ٷr����Y�RF�����E�6�\u����q��&�*!qל��~���	�'�~d�_r�M�ۋ���G�yn�N�N���\\2�}�0Q2��ݪ��_�'=*ڵ~<wh�AAu���������V+��~���5��_�5wn?踂��	q�Ύ�77���������c��7?�<_�|TxT��Y�[�V�T	+��;���:P�֮��a��m��IC�l�lb��?�-Z䒲��T�X��56�*H┲�:h��[��^��ör�/ʥp�X�n�[�ei�/E����V;�	J��e���鸩���yϷMM�۬�����,�t���#ҲP����
M���;n���M���V�g$��>�g�H^��7[-�Sw���ܡ���e����v����*��xr�M�wy��{�j~}o�]� ܬ�K��m��T���Eb�إ;/s��b��3k!Vj[��WV�
�[�j��vt�_w�/����FY���'�C�nO�J�|�7-ۈ��9U�#�7&�Z�02������l�en�C�$d�)m$�Ej)�<�f+!r�7+n#�B���?ݍ�է]��H��^g���۲����#���ɣ��+����v�������~H_-���O�V3rO��Ҭly1-(nwV���v�J�����ͣ'�_���s�6���V��٨ڵ}�W��j
�LL;V����qq��9}*��W�9{��7``q��/�5٨����5�;Y�Ս����^��7�^�ڷo���5ٮ�vk�]���f�5ٮ�vk�]���f���;��w�zw�&��ޝ�ޝ�ޝ�޻v�F�������|�͛5۷@��v��4h�  Ns��9�s��9�s��9����D]�V^դ���N��&���a�F�<9��Ϊ�֧9y9����G�$l�"���_��Ma�Β�Y��,���"����������\Wƴahï���R���V���ȥ�t�j��U���nn�&L�_ɓ&�F�ӽq�*?�J�9���ך2֍{;�t��Opդ�c�-)��r����F�����J���~n9��\F}�iJ�Qx���J�6�JUa��澓�lHJ�H��M�ov6���Ż���I���J��'F�ɓ_V�5gF������     &���ջF���L�2dɯ�:5nѫu2d�h�;ɭc�IcaI	�������ؽ�T�ݚk�o�ϝ}}}���LLM�V�ѣ}٦�ǅ6|�P��,�}((L\����3s��'��g�J�5�]��zY�l�W���}`y�����������D�K?��U��}����4����q?���$�dBB�n�%W(ombR�g�ڸ���֭c�W�\a���F��4U���V��[^|愁���8x��I�YaqW��|������m�4@���xsZ�q�5���l٪�k��X�JIV娙T&n/[M�I�,�MY�bm�W�+��9�nIJ��.V]F��\{j9�cS��#�,�2��lb��/���奼�3݉���f�[�P�{ڌ7Yn�l�9{o�复l��ۭ��a��n��/�҈l�7d)?��X�ʢ��C�r����lC;#B�՜�^�)ok��KQ
����gۦ�ҭ�d�1�f!��[vQ�/v�m�GemF��(}צܥL���e�V<���n��M$J���n��J���8�Z��4��j����"�۩�����w��"��*֬�L�Sv��o����ܗW)�N���v9��ě���Y�"ߔ"�>B��Yv9���/��J�w�N�B`B���$[����;���]���j��J��rom>=�(|���J/��H["˴�wm�)U-Ir�?��Q�te+)���V6�rlr�H��F������MyE�%H[7V���o�۴�z"��������p�Vݔv�����5�ܵf�l�l�2�_�����?~�u���3�=y����󗁁�׭�*��j23̚MI׭���<����/Ϝ�>r�z��׭�x��˰�=y��/Vw͛\2�ջ~�tc�q�6kXpգvk�]���f�5ٮ�vk�]���f�5ٮ�}��vwݜ�N��&M;ӽ;ӽ;ӽ;ӽ///v���wnݗ���V��0 nݣF���   '9�s��9�s��9�iΎ;I�.�v�U��;�ѵ��f�4�Q�;�K棢n���z�/9��Kݱ�I��Y��z�a������4S����_�]���A4U��78�,p_�,��lcz���~]ܖ�i��r�qn��`¤�nR��4�3@�K�Ǉ5�ɓ.�2k�o�/E2hO7z�ޙ32�7�:�,���_�������@��Fڌ�Ոp�;��ĕ)WʰS&����I�2
3E�M'�Ic��"�F`H�ݚ��(�d�? �s�M�l6����@��<�����ڗM;ٴc�F��΍[�mK՗�;ӽV^�     �]�|���jݣ|�&M/���7�L�w�&M;ɓ@�뫯�ɿ�ٻ���Oaɿ���fюw�h�	��ƒ��7kWݝYz7Ѣ ��I�YKsw=�z�I���}�_ac�g&�@��h�	撒2M&����cccg*��Y�P#����dj�B}��
�XO���1�Q�I��Wn���JR.+oZL	W��"�m:󵎮nr���Ǣ�>��󗄄��E^�ms�/�l���?Y�"����F}�		�Ϝ�|���7[R����}�xpڗ�jլ8��Ǉ��	d�Wn���q[u0���-Y�lm�[/ʧ@�S�9�)e��{4N�nW'ʒ){�,�v����iy�治�e��u�͍O�����]gk��~���w�*[��"�)J��!e�-�r���א~T�������d����s%�
�X���ZΕcc�e�dV6:�w�J����Z��+L���1x����òP���F���ZfK�C��[x�FD_c��PePݦ��[N�Kx1}��!�����Ӷ2��������Δ��c�vSw��-EvR��;�\�/���^ߎ�]>E��b����)S�qyM�*�cì��%Xp�6�o%���_n�)��d�1��K{��uψU�ݸ�o����ub�d��#{.,w7aRT6B��k�!,x�lK��nV�]���؟���7$-�v����V6x4�d������ވ͹*v��N�䐷l�:n��X�S�����۽��b�mo;��d�{
UJ!)oV�vU�u�9��_�ݦZF�|��(����ߠFɰ<��ǚ_�m������=l, �l~�AuѢ�Z�x�������s�/�E\٨��G6j9�QѢ�>r�|游Ï�yu�����������ю��8O00�`a<�ݚ��f�5ٮ�vk�]���f�5ٮ�vk�_vwݝ�g;ӽ;ɓN��N��N��N�� *ի�4h� �}۷g9�  	�s��9�s��9�s�sM��o0+��Q�Wݺ�5��{���v��_4\�Q?�c��2��R�t}���{#d���|�hNl5p��](�K���.��x�	6!w�4�������`«}-�ț
K�O8��
��N��pջF��΍[��\y�kF>��K+�4��t�<´�c�(HWe%rUX��r�;�����qn����]5�L��l��V|�3ZhƸ�'��'�����B�l0p*��'��g�N^��nɤR�y�a�/qךd�ݜ��h�F��6��ڗ�F�޻F�     �΍[�mK�/F���L�w�&��o�V��7���7՗��5Yz5�{V�}�R�Q?p0l��h���O,��j^���u碬�ɰڗÏq���D���maL�F63#�ss���gܸ�p,�p,�8xc�����{8xw;b
ݖM���+���ݹ@�����u��'�L�̟_�f��
���U�?dU��[��+Nw/��q�^��q���^��lo�<�3��82{��zȤ�-��.̋���]tK�f�Ϝ�>����qq��������6=��a��&�w���jh/lC��i�ial�K�.^=�N�ӷ�X���F��Jۭ��
����ӱ2����B�o�ɖ����W8����^O�UM�V7�����l���׶�\`B��P�O������}�G�&J���i���B���Y{���*�!{j6ݜ�N���-�Y������vW�C����n�v?�υr�I���g^?����v�R7��n9e|+o���k"���[)�eퟒV������2ؚ�R���QX)�liY-�z�ݡ�ӱ14VR���RD��[��W�����o*��Tpi�yUc�(Vt���JF�m-�}��ݮ񳵚��#D4�~C{'ېy��W�.�.��V>B`\�/{�Ê�r�7�/_���ry�\����&Fk-���J�E{+9+�l��-ڴ�7�!�Yr��������i���J�G��0���g-�i�̶^�q�b�IB�Vۚ�u�Ow̙��E���V�$ߘ��zv�H���9�4ܶ��?T��i)!>����/��n|��f�qq���|�ǎ���f���V�Æxp�ի�㻛5�n>����63�k�lv��F㝯�=a<���sюթz���ݚ��f�5ٮ�vk�]���f�5ٮ�vk�_vwݝ�g;ӽ;ɓN��N��N��N��U�Vs�����>r���9��۠  ��9�s��9�s��4��~������L�v^ա�5�6���ݻ5�_4��9{�͆��Kѻ�F:5n�Q��㝮�2�y}162�U�X�F�j��^�ש0$�[w()=z����R��-�{
:-�������2��o��&�ǆ��ɪ�ѵ�Ǟ��n"l),$R�Ie~���&ͯ,�۫qɑ�>��r�B��$��N#n�m�"�D�ٳZKն�d6��Ź���_��"�`qn�RF/f��W�Yf~F�&��O10V)4e%%�}�O�w*�ѝ��΍[�mK���##b`|����f�2i�s��9�s��9�s��0'9ݻv�۷�|�1V^��hջv��ݜ�&MF��6��y5Yz7ݚdɩ,cll)&ͣLddlJk�o�	�Y&��F�՗�������V�kXe�վ��'/�EXɮ���226E"�I_��"�J�W)gd$�O�X�I[M�#c����NW�/��Uz��a,�G��p���KsnE����{"%;;,�X�P4X���j��P%Z���旫8���qݗ�|���f�׭�HNq10110110?�����t�>c>���V���q��
�Lo����b``|��q�������Rs����'_�����[:��F��;H��O��l�-��߶=�����\V!��gd�=�e,��ȡ[,rkn}�a�Ev�#�R�o�)�U3k$A�?lSǐ~QO̵+"������!�K8�[%���᤹m�;�7v�e�S��Y"!e�nE�{�}������Pܵ>3vP�����2�nvH���ɢ�H��;�[�ju��NDCeX�۴��*��!%e8��	K�lҶ�y���{1x4�7-O��(4�w+�␾\R�nB�v���]nnK�*���v7��&�%��%mGV����k��YQ����W���~>/����L�Sݯe��659*��2�	*F�B���:�����K�������,�̖�J�V?*�09$+��Z,w%\2����I��qSd�*��7%�6:��R�|�-r�l���o���D6�WiO�R�~���?%��j��P[���Ƶ�Hњ��;[���e-mNە��P4�4�X1��Lv&�*v�� �.���5i҆»�N�XnE�-�^O�r���L�㝭��ͣZ�V����ׯ[Wn��F�6j5j��F�6j=zڸ�Û5V���h�WF���|��Q������g����Y_aV�����n�FԽ\ְ��kF;Z1��k��n�vk�����xe��ݼ���5��ٮ�vk�]���f�4�9�s��9�s��9�s���9�s��0       Mag"����cH�0jݣV�[��_5�Q��/|���F��vwݚ��F��oU�<v������$lL��D�^^U�FpU��k�0����F��i2l0=n ��ɫ�75��3&��씴�^;-�K��d�e���½I_c��<9�Q�V��}�E:�!�r���ȉ�n�bỸ�l��v�VU��N皯��~�XIe~o08Y�2)2��Z\<��f[g��D,����z�������I��f�k���h�q�kTj�L�5�gF��=y�h���7�L�w�9�s��9�s��9�s���;ﾍ4hѻv��1}����N�dɓ&L�4���jݣ~<ֻ7u���.:�M_'��������/E5�n:��	�G<Ӽ������5�k���Z���'}��M���"by(��:A��݁������ݕ\�[���ol����|�T�B�!P$^���K�r�V�+��]GM��/M�6���/S�
��G�.+n�BP��v�[F����/~/>sD�������54V�_���&�<tsa���xH�|����j�n-����Np?�u���_?�"l"i,��8���Q!��W/]�H;:U;g]�ji�Tܽ�+e�o���m-�ĕY��ȭ���w�YKL�}�a�!e?����v"F�er��O���\�k�
�R�`Ӱb��/��M���^��+Q����D?�"��m�-n���FJ�w*w����g�6����Ī�cɈ┱2�n���-Ö�JX�/�V���"���D$���-�V~$lW�-��E3���3��b����)/ʥ"y%V��d����I�4���+Mg��ᔶ��n�*��9%,�+M#ji�=�*�좶}��]3SY�J�����p|F^�F3�>/�ϋ�b������X���e���۔7M��)W���Q}N��O�c�����c��X�i���#Q,��[u��l�-��Z��%ldn���O�F?�B�J�V'��[�ӵ��fε���~4BJ�e�pL��������q��T5g���2���_#�M,������n����Rk�$�v��F��)wmI��.X��Ε���p�|G�����ҹo������^z:�c��:�X�݁����l٨��GϜ�~����[\����Fի���23̞O�5*����Fy͎��7W�/Vw�y��ְ�Q�}y�|�ݾ���ݾ�󼼼��v����yyyyyF��^^^]��חf�5ٮ�vk�]��Ӝ�9�s��9�s��9�w�|�9�s��      |����K �,m\sQ��7ݣ}[�Ѿwo_5��oK�<7�^���:7΍���;�ݝ�oQ�}�4y����X�H���~xq��w5Yګw6�=t\D�_�z."`��sL��&
6M^�;U|��N�T���݇�-��J������4�<+��n.�ѫj^_|xP��e��s_"�����һ�X�q���D�.N_6�i�wv �<5���*&�����������4�dR���`jᵎ�i�wf������|�ݾ����yyyyV���n�s��9�s��9�s��9�}�nݣF�4hѣ}��s	�&L�2dֱᵏ�&�j^_[X��������ϕ@��Խ��&����MV^��xnѽ2k�����EF��חݝYz8q��Ϟn�9���X��%�ryV�B����Y�ͻ=���b!HY]��B�e�77,%ZR�.M6ϻ���y"��)e��Kw"��_��g�k��������S�,�w^e�G�QyKi[�wd6�w�?j�ȵ��]�oa�;�pQ�a ���/j��4U��4dg�x��j��5_�tF}��������}�q�����������0PP]|����&�Ug��s�݄����oy!z+�-DJ���2ԫ�T&�K�J�i�o��^���)Cu4�8��Oô����b�Lv����[e7[Q�����'�hw����7�Z��*�r��b��/[n��6�8�Uc̞'ݐ�\RV�w�P�����߶Oé�lb��~�o+Lא���W�;OϏ��)ފn�[Ϗ��I��Y.�fR��(��\��7{S�e��t�_�J�e���엒�0yJ��Րu�\M3�����u���M�p�X���_�%dV68ݤfܕ���J��7g]�o�i;%
�)*��P�JZ��v+�N��q6��Nt��[�����{q�W�Y�a�� O�4�[�����Y�M��lwkx�^+.�U@�f�o�϶�yYI?d~�#�n���$��J!����rW�*AX�Yw�,�;���wQC����b!Y\O����QZ�*��X�@�B��}5f!%j"�lM;-Y��6ܯʛ���ܤ�ݒ#��G���7i@��|��e�2�l�ݰՈk��._�zI<�5��tf��3������8gϜ��MI��_�������իWժ��^��'WW;��Q����6:�h��_5�_5����<2�z�u�����;Z3K��v����/Vuh��]�|��v�������7΍�5ٮ�vk�]���f�4�9�s��9�s��9�s���9�s��0       ��U����2&2���^��u9�vs�;�ݝ��Vw�_4����^wѾto��g}��V��޻5�n�͇<������cq����f�wcʀR�7{xWoM"�����Z�ܮ�Y�
����8�JL	6�HҌ��З����5�j�MkF??�bc ��~��j�`m`F��Ƞ�%P8Mo�Ϭ��o�E��V����RX�H�����II&�XʥV2�U��ߛ6}��ca�����e��G�������V���n�ѻ/F�[��^^^^]����գ9�s��9�s��9�s��v�۷nݻv���9�ɓ&������Ѿ_[�oL�2k���$��Q?y�h�V��S&���K᫆Ժd�ݝYz3�/Vxe�/WF;Z9���6x���_"������)ew!��-��ۯ��P#�	A�V8k�~�����89��K+���䭖�sn^�2��U�a*ձ�������8J��BM�\��_���k;ܝ��M��
ue�浛[UXj��������AAu��6l�pᝫW�f�	�6
6
�<���BXF�������8���<�0������_4��}\��b%z%.�!oe�{-���ܥ��b���v���۸d�eS�壼T��&����ba��M+�+Z�b�;*����vQ���Cխ� s齒�;���TX�H���j�ݮ��rqFOݷ�54��/ɣF��?��JU�x��[O�C�M��u��C��TduYJא��ZԚ��P69}��;��Y@�X�����~v�)���c�wY��e��R��8�,L��z(~>����-�;/ �)�Y[��7�}��%Va����%��[v��cco������JFȧo^t���f��B.�@ɸlt��P��ӋXv)�u�-+m$��)n�x2Z9X��xc�L�L��^˷X����ͺv�n����(|���eQ{V8d�0�������W�ė�4�mE;-Y�Su�]��R��x����
E@���D�����yJ���d���?r���ܲ��6��ݔ�nPߐ��������dB�Q9�	T*B��r��vH�&��a�/I��[Ϗ�X��䃱�D$�nW{��;b�~�߿qᗗ�w���վ�l�n.0��/�E"�������$'?>sh�V�U۬x��Au�K#p�Z�٨��V���њ_6:�oh�/�6:7��^��z7o!?�B��矘�f�V���gk�2��՝Z*�R�g�^�2�ջ}�����vk˳]���f�5ٮ�vi�s��9�s��9�s��;�s��9�`       ���7>bb����9{V�պ�2i޾^wh�z��Ѿ�y�F���:7������vto]���F�[�pջj_�%ě"E��K%Ro����V[g���*<��8/��]ћ_�4�z���^�H�5z��<p�7贫z�^�Hϰ1�n ���jr�S_vr�j�᫟@�Rn`�ғ�o�`E��.Y��~�ڂ�I�4�p�����݅B�uu�s��	Ic���~ո��__���'�����IcF�2d�ޝ��Q���o�V��z�jѫv��^^^^^^]���|�9�s��9�s��9�s��9�s  N��g}�ݣ}�j�ѫ/Fw�ջ�Կ�O66�`� �~��dy��5�ɥ�ի/E2d��j�.�4���j��矛�|�a��k��X����ǎ����k�Yr����m~F����WrP�쳻��F��^^
Yg
��dZ��n<�D"�;�r�-������M����
�g�z���o�v����ġ��l69zַQ$m=�.��5p��qV����Y�Q��teֳQ��7�9��}��a�?7�`�k�>�D������y����7>r���Î�\�?a>���7XH�f�~�e��8�K�Q�죹�d�ݹJ��*�[�����Wl�YՋ���O��\�.+n�B���[����G�R܅��d>6Ε���e����ҧwnR�f�ݠ�Z�t����R�+;Z��9C�Q䔲��!��1�=�����e�R�-���C'�a~;��l"��!������r�-5&�v�(H۶\L��`P62��d��M��q(�f䕯 �$/l{o%#uϐa��en�7e������S�,��ͥ'R��_�!l!����v���R�Z�����V��
��Pef//��V�nRUŜCYY�k��-n*�*�ʑ�2!�d�p�����F��;3��+l��Q�:�D5��d���f��ېv���(oj6ݔw�Eo�Y��%����ҧwk�4�Ȇ���K6�,1�����x�.r��"�f����m���F�Y�
�P%��C-'լI�+r+���bub�Q�)�������r�϶Pᔵ�r�^���܋�n�,.V�k�L����%g
���*e;b�E~2ʹ���&�H�ccsK՗�����Th�h������\\a͚�dg�v�_V���GF���QÆuj�h�Ϝ���h�9�����<�ڗ�F��F��EV�^����^���]�|ٱ��j�;Tma�k�v���WFi~����/�����^���:%��f�5Y��Vj�]�s��9�s��9�s��9����9�s�       9�s�8�����8j��2e�������7�}��}��}��}�ݣ}�7�vwݝ�f�;��to^�a����Ȃ�����h����}�O��Y�Vrr���_�qn�`H��%V{t����ɫ�����}%��Tf�w�;�ϲ�<�h�Myyy�e���X3M�3rU	�,u̗�c��,��s̽�Y,�O���y����������K%[��2i�Uca��ڲ�n՗�V���_/;��}�V��o�ٯ//.�vk�]��ח����9�s��9�s��9�` ��v�۴o�F��o�V��j�ѫ/F��5n��Icٻ�ɿ�&�K##beY?�<���L��[�e��vue覣V��e�՗�k|5o�<	5�$O�z0��w6��<����I�&2�Y&�G�����:��2��C;���(jvT�*J��Ȟ�\���^KDiw$O�	f�*/@�e���'�Eˇ͆��4��O�����3��L����Ci���m�~���L8���k��o��=e����7��a9��k6j9�QѢ�>r�z����:>���Ώ�t}��YᢣE/.���_9�"���}���������e��e.�A��xr�K�*3oc�%[yT���)�(Vwc��V�v!!l;!Y�Ig��4+^/���e��C��I�����P�EP��i�ڜ+;Z����/lz۱�ӻ��j�)Vc�Kn��g��Cv��,M�iJ��i��+''�exqx�v)ܹ�����r��]�Qە�~i���d���Ե��t� �������i���Q�%S!��ʐ��K|��{tժv�����n�;.�)���d�~�vC�[�v&��b2�]Mk����,�(V�F��V{r�=d��T�R�_�����$��*R��P2���'S�z-�<�[��w%�Q8�l8��i�2���/(|����n��%j!�_E%�۔�|�VS^��䒲��&��R��!��nJ�8n�E�`�3�Y�zƦ�� ȸq]�O�;���ҨV�!)Vu����C-ken?��~H?-Ⱦ�O�(c��Z�`��U����l�,x�w+��Y��*4O�^�ϒ�/��n�s�*n��|7^���I:vZ��!kz��J?��������"a ��a�;�U�Æth��^��)!?�ћ5x���/Ϝ�3���y󗌌�cc���<����V��c�G{��7�^����k�k��޻z��v��F�����j�lutf��'[���旫j��7o��tJ%Y��Vj�U���f�5��s��9�s��9�s��}��s��9�       4jժ<x���GZ8j�V�e����诽}��}��}��}��}��;�ݝ�g}��vs�;��tK���=q�N�X�e���g�[�{��6\FVˈ���mj���Xj��i���j鎭o���2]����0�){���ݷw�~�Ug����c�//F�<2�p)%�z����gc�,��D��1�4Q�����7o�ac'�����V_4��l^�!b���&L�2r�jᾍ�������ח�����f�5٨�;�^^^Ns��9�s��9�s��9�s Ns�F�8q��F��5nѫv��Ѿ�����4ӽ�ԼLdm$e�S���Y&��D���ɧ{�Ɗ��gzw����j^����pڗ��W�D��lu`|�����H�R��TC���>�^[eN����ie��c�#?o�2���66O'����c'.���^Y���m��e�bR�o��y.�݅j��ls�#�-��~?����N^�&ue��ǛF;Xn�G�\q�\�bn4h�ϭ��su��9�!9�Au�������]tK����ΈϽy�j���c�v�����HȘ��ް?d�m��"����r�N�g۳ϭ�u��T_�
�S)���ˉ���H���/�����Bvu��dv�-���o[��-��3r����jnX�on"��M�p�$�����*9�/'������|+S!�"�w#T����o$уIr�0"�v���{�ǃ(äw�;����l�ߛ.��'^���~l��:�6R��E2X�}cg�Ȧ�ϐi�ڝcg��w9/ �S���W��J����,�3^P��==lW9�[���v����t�7�#v����e�$�$����ga3�Q�W䥰��P091y�mwQ-�{l�ۉ?$��*��$�_-�!ocw+y�����P�@��hxpi��辶���~���uo��+?Ȇ�
啯��qd�n�����}�/���)e�a��l���V����NB�G��n��J�?�H98�s#�9Fە���ό�~j��Rm\]~�._��}n���e彬1���w���N�*�������f�s����[~/g$dB�(�(��,ߔ=��C��!kv�
V�%���M_Iacc�
E'����q		���3�E��.0����9�.0��W;��_/.�EϜ���JHJ���0:9��q��{��yyy/F�z��v��z��/~{��߆^�z���:�Uh������Q͎����a�F���~�՚�Vj�U���f�5Y��vs��9�s��9�s��9�}��9�s       
7�vs�v�7g;��l٣##/�w<������/5��[���������}��_zdӽ}�Ѻ�uv��]�EU��;P9�d�9��c`��f��J���U���s�W�~E��c����2%b�����BW�g���W�g�ʤW����3Dg�7f�G'�5|���ӽyyve�+�1�^qڌ��I���П�n�K+�������w3s���e%��m����$Ш���/�E�6�ᵆ^�Z2����/j�uS�Q���^^^^Q�to����ٮ�yyy9�s��9�s��9�s��}��}���4hڵkF�z��F��7ݻv����&Ç�7�X����to�Ϟ��gg���%}���_}\8h����W6�i�]�|��ݝ�ts���;������������J��px��i��[���*�6�!�_�nˇW�W�ϳ����v�I���)e�B/��lm�\��*/��{8b�z�Q
n�/O���gv�S��j�AF��[���|��j^^��z0���^tn4]�����^�*�g�����?��͚�%$$lo��(�ty���D���P�9��>�Bs�����k�i5%��L$$Lf��ldڼ6�E�J��tؘ�Kr��i�Jf�;��2��NF�#����5��J��r	8�1:�:���[���ᒵeQyT+M_�(h�B���-�/���B�Q]Y
F�z ��1!bn{�kv��#iJ�U�Q� �*���������;9��d�������!YY"J�ò����vݷ(H�}�ZH��v5؆�����qb��lWVA�V��8�L��a��E$���M$mrYH<�L��9V�v�+�Hp�L��S�ܧ��Y{�1셽��2�������!l�ܗ����r�4�R)�6-���ci�S�t�����%��od8nʵ"��d�CS$S�V�U�Q���)��}oas��b��*����ϲ�,;y\:h�K'R쐲q7-6��M�G���vB�P�qN����6��Z��L�'~7_��������d��7en����岻:�Z��f�n����|;{�In�S���rdCdM؄���ob�nA����V#a���-��=�@��s���SX�{i҆�?~2��O'���J�r4�e�|�o玍���<�3Ϝ�4U���
�>r��Q��^���W�z��h�f��5V������kV�͚��N�~�]�V����Q��;�^Q�w�v���R�gV������޾k�z���j��/V��f�4���v�{�Vj�U���f�5Y��vk���9�s��9�s��9����9�s�       f�j���F���Ns�����p7��0V1��4.��f�z�뷯�}��_}�ޙ4�_vuh��Q���R^p��z�@����������W����Ƒ�]6��i."`�[{���l�t]��	�,@���Ջ�?9;!���_��8a lr0 ��'F�6��s͏5�l�ٯ��DLLnL�Y"�D-��^+��~�M��Ea"�\@����<q1165���03�t';�s�����vs��T�U;�        	�r���n��󯯯������Ï��q���<d����D������^b`�Y16��3&�/:���ѫ/~lun9�њ^��9yyz4hݣ߿e��f���}}>|�77!��oe�o?�v�Yg9|k������C{;h��,�WrE��'��a�k�N��7��gv��m����n�g��xk)U��lkV�������	_��ő���Ǟ�z�u������n�2�z�����[Y�Q�j�V�Ѣ�$h�K��q����D�<tn1с�/������c.#l?�,�ll?������OI	�K�nU��,��׈J�4����+�7w�ˈ�d��_��cg�	I���?9n2#0!���_�!�M|$��^?�@ʳK.�ȸ���'�D57,^NE��e��T������/����<�$Rᾊ�A�ʲRD��݁����;����Ǔ��A���8�h\w�S������aR��H�p%��/���d�p�U�eJ�J��7�M��z�#⁖�o�}�knv�M�Kv�U+eJ�ge�b���Jz�����nL�O�n��X�C-O��;d��+��r��z+6_6^Գ�4��E�e��2}�]����ӵ5�>����V�|�D�������]f��|k)�zn��r�}U�!����uVZ�Eo'"��x�Q��^S���"��~+e�G�4�b?����m�4�v�K�{�����!�>χ-�M���
���Ce,�fE�������ƚF�i��)X�Hv��ی�o�Xmw�#���c��8���BO��|�E���;r�v�RW�>B������O+���Ӷ[��R�l�V%�M~��U���z(�A|�^Ug��'���qq���>sD����q�E^|������kV���f�G6j:3Kբ��Ç����ՓRRBB}ͣE[V��UV���w���gv�Z,2���v��e�v��U�}[�Ѿto��vk��٨�:�o�v��o��v^��z7e���V���o�ٮ�vj7΍�5ٮ�vk�]���f�|��vk�^^^^      9��F^�z4e�Ѽ�F�<x�s盟<<�a�<ӻvto���5nѫv��z��o�٧y4�_vwh�}[��]�[R������q�5����ڗ�q���^��a"~���$�)e��O/�G8/��1����Ay�'���E'��"�����nvp����V�e�m���֌�%�R�?���1�0�2}�7�dY��V2�5�� �y���V��V�9��������v���v�����vs�9ݜ�U:�ݜ�         (ѣjժ�jݻwF�������a>�ǚ�Y|z9����^�2w��9{X�V_���i,h��q��M,����\�>y���	j�v��V^����ã4�����ի�6o�~������ȤR(HHL8p�iidij�$Vv2�7���8������m��-l8�U����䛲�W���62̍{����|�JE���@���-����g�����)C���vR��u&'?�x(�=~������`n9��u����2�~������th�׭�/��`������]����VD���_�p��k�Nh��?cy��F�;�η��z�
n#-�r�5��}�X66���
�f�$m�;��w�ZVnD~ϲ��e�g�i��d�7$�	�
�&�φɷi�R/ϲn��}����Y�L��BMm�JYM�f��쥿�n�H�ok�2��ԡ�:^~V�_�iHX�n��ŕ��V�1��8���z}u
P�[�W)B���H[�nR�PaYjd�������i�rA��ϧY��)��?$�I�M�p�d-dv!(e�x�Y�@��u�_�vF�li�*ƶ����gi�]������n��({b��=���!�8��//�)bl�)7��7^O�X�φ��UK���h{���۴Ȑ��P��&����aZ�T���;+tC+Y��(8�D;�Y]��Wv�޼�Z��0ݕN���b�6ݕ�"�ݲ�`�糮�K|���0}����(<�D��c�l�&J��[_ud[���{!��JeK�G;[g�%`²�rUf3vM��쐵���WYI&�h�a�&���߰Ȉj¥-z�wW%���l.R��nR��Yxl����b�[�g����`�E���*�k��z4lc!,c?�\a��4dg���y��ۏ>s����P]bb`a!9�����9��u��k�ۍ*�D��ҖF�@��kG;���˪˰ᝫWᗾ^��ޫE�^�Xn��w��n�vj�o�v�7΍�}�g;���΍�|�ݾ���ݾ^��z7e���V���o�ٮ�vj7΍�5ٮ�vk�]���f�|��vk�^^^^       /���n�ѣ/F��7��j�͛7>�n `s@��q�to��ڲ�j�ѣV��7Ѿwf�|��9�M;�ݜ��}[�jݾ��ջ��n�7�c�/F���ݝ�7�vtj�ǚ֎y��/j������idҕ}�ױ�۱������JU,������I�����V�=
7���'쾌r�.���<�J2�7�*��m\u��Y��c`��|5p�h�p�jԼ����}����իVs�����vs�9�N�uS�9�        s�<x���jլ8p�͚���|�Ï6y� |��q|wf���n |����Y&��`��q���+L}y���M*���������%5h՞l7��/�F��ݻv�Z�jկ���P(���PPY�f����J�Q�6Q��`�ms����M*ҏ�e.W;�2Y!i����{m���	%��ȹp���XI�ViW8�6F䅒�r�T�CS���rXg�d����f���K���J5qݣ|�O��`|������??�B���ǟ9�`q��㄄�c��\~n-u�/q��\�`tK�����wsu��XL:1��\q��n9������V��ܶ�C���#$W/�X?�ɮ l%�AQ��jH(�|(���Kn������rI[���+%�퐷���l+���v�ݎ�_-�ɋ�"�H�qR'>A���Z���Y�vul�x�/͝v���o�cЭ�sMn�b+R��ŕ��8�S8����/9�qZ�Ӭb+8;�T+%�ն�i�<�*���r�딡��X���ɷ�ݖ|_Y_�!Y��Y���(lf|��N��edi*������B�ݒv��%� ���;nP�ܱy<�&�!{c�:엔�j��S��M�K'���p��+bunU��#�A�YurT�����-��ca�{a���Tn�"M���m�8�
�;e�E"�:o���������;|����9���$8˖W�R�B�Q]LvK�)R_O���u�(M)�s�M����/��ܐi%P�M(����"�)e�\�T��Pېw��I+ML�l��Ԫ�����_)"�����ck�6�w�2˕�cw��z-�T���-؆[��r��N��Ѵ�m��.�P�qP"k����j��Z�j��P]e���(.�08���׭���(.����b`l, ���cc�Au�I�"`�������Le�F|�
'��Z�9ݵ�V]V]��Z����gv�Z,2���v��e�v��U�}[�Ѿto��9ݜ��to��F�ջ}[��ѻ/F��jї�v��5ٮ�F�Ѿwf�5ٮ�vk�]���o�ٮ�vk����      �:�n�ѣ/F��o/8`��q	���;��n�ї�V_Y|5j�ѫv��o�v�7�w�zw�yvs�~R�ݜ�U���Խ�o�;�oMF��5n�MF��5n���2j07��?���n[+Ý��1t��+r�X�ϕBH���if?�mu�_5[��W5�}�