3480
700
700
3
255 1
1 01
83 001111111
74 001111110
131 001111101
175 0011111001
4 0011111000
37 00111101
209 001111001
166 001111000
0 001110
58 00110111
127 001101101
22 00110110011
5 00110110010
172 00110110001
55 001101100001
107 0011011000001
119 0011011000000
220 001101011
194 001101010
151 00110100
101 0011001111111
120 0011001111110
128 001100111110111
138 001100111110110
80 00110011111010
86 0011001111100
38 001100111101
133 0011001111001
104 0011001111000
2 00110011101
66 001100111001
17 001100111000
19 0011001101
147 00110011001
105 00110011000111
146 00110011000110
70 0011001100010
230 0011001100001
150 00110011000001
181 00110011000000
240 0011001011
92 00110010101
42 001100101001
106 001100101000111
82 001100101000110
130 00110010100010
102 0011001010000
12 00110010011
23 00110010010
97 0011001000111
64 0011001000110
144 001100100010
180 00110010000
108 00110001
207 00110000
218 0010111111111
85 0010111111110
116 001011111110
20 00101111110
223 0010111110
50 00101111011
179 00101111010
94 001011110011
202 0010111100101
81 00101111001001
125 00101111001000
41 00101111000
243 00101110
67 0010110
117 00101011
32 00101010111
118 001010101101
62 001010101100
34 00101010101
221 0010101010011
142 0010101010010
65 001010101000
51 001010100111
49 001010100110
155 00101010010
3 0010101000
182 00101001
228 001010001
195 001010000
244 0010011
69 00100101
232 001001001
239 001001000
24 00100011111
152 00100011110
168 001000111011
198 0010001110101
76 0010001110100
139 00100011100
7 0010001101
31 00100011001
54 001000110001
45 001000110000
254 00100010
99 0010000
60 000111
234 0001101
8 000110011111
84 0001100111101
159 0001100111100
16 00011001110
48 00011001101
25 00011001100
171 0001100101111
143 00011001011101
190 000110010111001
95 000110010111000
46 000110010110
124 00011001010
13 00011001001
73 000110010001
187 0001100100001
112 00011001000001
205 00011001000000
236 00011000
153 0001011
68 00010101111111
241 000101011111101
178 000101011111100
154 00010101111101
186 00010101111100
30 000101011110
63 000101011101
165 0001010111001
129 0001010111000
224 0001010110
136 000101010111
88 00010101011011
122 00010101011010
57 00010101011001
79 00010101011000
163 00010101010
15 0001010100
18 00010100111
229 000101001101
191 00010100110011
162 00010100110010
145 0001010011000
204 0001010010
188 000101000
247 0001001
44 00010001
199 00010000111
35 00010000110
208 0001000010
36 0001000001
39 00010000001
149 000100000001
110 000100000000
200 000011
53 0000101
135 000010011111
78 000010011110
14 00001001110
28 0000100110
6 0000100101
183 000010010011
174 00001001001011
61 00001001001010
113 0000100100100
215 00001001000
248 00001000
9 000001111
216 0000011101
27 0000011100
29 00000110
11 000001011
211 000001010
196 00000100111
21 000001001101
109 00000100110011
185 00000100110010
192 0000010011000
72 0000010010
176 000001000111
75 000001000110
114 00000100010111
156 00000100010110
177 0000010001010
167 000001000100
141 000001000011
160 000001000010
132 0000010000011
71 0000010000010
87 000001000000
52 0000001111
59 00000011101
33 00000011100
91 000000110111
77 000000110110
184 000000110101
121 000000110100
115 0000001100111
140 0000001100110
170 0000001100101
214 0000001100100
103 00000011000
47 00000010
10 000000011
231 000000010
43 0000000011
40 00000000101
90 0000000010011
111 00000000100101
158 000000001001001
238 0000000010010001
237 0000000010010000
100 000000001000
56 0000000001
26 00000000001
93 00000000000
vinicius���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�?�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$O$ H��"B�$ H��"B�'�$O��	����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"B�$�2aD�&L�2dɓ&L�2dɓ&L�0�"B�$ H����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$H@�!D�	$I2dɓ&L�2dɓ&L�2dɓ&L�2dɓ&L�2dɓ&L�2aD�	$H@�!D��"�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$ H��"B�&L�2dɓ&L�2dɌ&L�2dɓ&L�2d��$ H��"���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�$I2d��&L�2dɓ&L�2A �$�@C�H```�H2��,�H2��A �2dɓ&L�@�!D�	$H@�?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"B�&L�2dɓ&e�d�������������������dɓ&L H��"B��D��"B�&L�2d�	$���� �e�	Y �e�&L H��"B�$ H�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$ H��"B�&L�2dɓ&e�d�A �$����I$000000H$dɓ&L�@�?����	$I2d��,�I	Y �e�&L�2aD�&L H��"B���	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$�2dɓ&L�2d��,�2c�H``````�$	�&$H@�?������D�&L�2c�H�II "dɓ&L�2dɓ&L�2d��'�	�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H�$H@�!D�&L�2dɓ$�A �$�@Cɓ&L�@�?���������&L�2d�	$�$�$�@CY �L�2dɓ&L�2aD�	��'�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'��"B�$�2dɓ&L�2d̲A ``````````````````�2aD�	����������@�!D�&L```�II "I$000000L�2dɓ&L�2aD�	$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H���&L�@�$ɓ&L�2dɓ&000000000I$��$���� �e�&L H��"������������2dɓ&000I$��$����������2dɓ&L�0�"B�$ H��"���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"B�$ H�dɓ&L�2dɓ$�@D�```�$�A �2aD�	��������������D�	L�1���I$I �  ����H$	Y2dɓ&L�0�"B��D�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2dɓ&L�2d�	$�$�$�@CY �L�0�"����������������D�&L�$	$�$�$�,�$fY �2dɓ$ H��"$ H����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�	$I2dɓ&L�2A �$����I$I$��	�&L�0�"B�������������������@�!D�&L```````````````�H2��,�2dɓ&L�@�!D��"��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	���D�	$I2dɓ&L�2A �$����I$I$��$�2dɓ&$H@�?���������������������&L� �e�	Y �e�&L�2dɓ$ H��"B�� H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ H��"B�$ H��"I�&L�2dɒ	Y�e�	$������� �e�&L H��"�����������&L�2fY �$H@�?���������D�	L�1���I$I$��	�&L�2dɓ&L H�$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��"x@�!D�	$I2dɓ&L�2dɌI !������dɓ&L H��"����������񁁀P(d�z*EH�"�T�L$���k5�&O�����������"I�&H$c�A�L�2dɓ&L�2dɓ$ H��"���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"B�$ H��"B�&L�2dɓ&L�1���������������dɓ&L�2�����������@�# �P(��dC.��bbb	@���x�����/��*EH��$�@AD�����������"I�&L�2A �$�@CY �L�2A �&L�@�!D�	������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O�D�	$H@�!D�&L�2dɓ$�A �$�A �$�dɄ	������������	I$��f�X�P(*EH�����~ �@����9NS�%�H�� <� G�
�Y�``c����������	$I2d��,```�II !���A �&L�2dɓ&$H@�!D�	$O$ H����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�	L�2dɓ&L�2d�A�000000000000000000L�2d�������������D�
��|P(
�R*E�_��~?�03L�46EA�9NS��9NP�|�`�!�1��~C(eblD#I$L�?���������$I2dɓ&000I$��$������� �e�&L�2dɓ$ H�$O����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"B�$�2dɓ$�A �$����I$000H$dɓ$ H��"���������� H�dɗ��bU
�T_��_���� �3$G̐,	A���r��)�r��)�r��(,	�`� M��d̙��@�Q(�I�&$O���������@�$ɓ&L� �e�I !���������,�$&L�2dɓ&L�@�!D�	$O�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�< H��"B�&L�@�$ɓ2̲A�e�	�,``````�I	Y �e�&L H�������������2d�0�8�B�����������0L�`���9NS��9NS��9NS��9NS��	A���f������2�Q�6&�BA2d������������D�&L�2c�H�I&L�2dɓ$ H��"x@�?����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$ H�dɓ&L�2dɓ2̲A �e�&L H��"�����������dɔJ%��U
��2�Q�2�T M�&	�`,��)�r��)�r��)�r��)�r��)�r��)�r��`��U���bbbfLə(
�D�2��������� H��"I�&000000I$��$�������2dɓ&L�2dɄ	$H@�?�	�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"B�$ H�dɓ&L�2d�A�H$c�H�Id�A2dɓ&$H@�?����������ɓ&Q(�CC�blH�#� @a	�`�6G)�r��)�r��)�r��(J>B>6eTT�1��͑�r��)�r��)�r��)�f��4f����8G�2�B@�������������D�&L�$	$����$�2��,�H&L�2dɓ&$H@�!D�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$ H��"I�&L�2dɒ	X�������������������H$&L H�������������2e�D
 ^��#�q�`�&��eA�9NS��9NS��9NS���͐��y�*����dU�! ���2�C"U�a4T#�0�|�)�r��)�r��)P| �`�YW*�d�b��_��*�P�1Q(�I�'�����������&L�2d�	$�$�$�@C�A�L�2dɄ	$H@�!D��"��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O� H��"B�&L�2dɓ&H$d�A�H$c�A�H$dɓ&L�@�?����������ɓ&000�� ��G� @� �L �3���r��)�r��)�r��)��π�#E8Ld�M�`�"��:h^fd����lDc`� #X�����R�zn38Ld�`�d#L��r��)�r��)�r���:d����4ʙS*G�
�Y��2aD����������dɓ&L�$	  $$�A �&L�2d��$ H��"�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O��$H@�!D�&L H�dɓ&L�H2ɓ&H$c�H`````````�2�ɓ$ H��"���������� H����t	@��8G�x,X� ��3LД|�)�r��)�r��)�r��6F̪��z88*ȫb��Z�����<����VR+)?�h���@�g�e'�BK`� ���*�@hȕr>g�8d�h<�9NS��9NS��9NS�Tp ��"�/��#�;AHR�������������2dɓ$�@C�A�L�2dɓ&L H��"B�'������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D��"B�$�2dɓ&L�2dɓ&H$d�A�000000000000000000L�0�"B��������������t$�I���3&d����~? `d�����t�9NS��9NS��9NS���͑�*����
A 	J�φy��$�V
�O�Z�=*�5�YI����VR+)?�����O�e'���A��̕A
�
OM�a�*��J>S��9NS��9NS����t&	�a��d̙�@�Pk5�ɓ'�����������$�2d�A�000000I$��	�,�2dɓ&L�@�!D��"'��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H�$O$ H�dɓ&L�2dɓ&L�������$�&L�2d�������������$H���:��@�PT��R/��/�����`�f��)�r��)�r��)�r��(<�3�0Y�6eTT�y�*b:PA �3�@�x	��3謤�VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����lD`@q��e�2��|�Fp�G�`�4Μ�)�r��)�r��)���0?���(e�blM��``I ����������$�2d�A�000000000000000L�2dɓ&L�2dɓ$ H��"x@�?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2dɓ&L�2d�	$�������$�$�@D�A�L�2dɄ	����������� H����Y��bU
�Tg�? �?�`f��h<�3�A�9NS��9NS��9NS�F���#E8Ld����!�*���g�<��(�6"1YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?����H|��lDb�3%PGB��23A4S��L%�)�r��)�r��)�T 0X,d��� @a `�H�"�@�_±2d����������@�!D�&L�H2�	�,�2dɓ&L�@�!D�	$O� H�$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�	$H@�!D�&L�2dɓ&L�2d�	$�$�$�@D�H�I&L H��"�����������L�0t	vG`�2�P�?����">d�`�Y�r��)�r��)�r��)��!P�������#�U,g��3�@�e����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?����A	,U�(�3�@�c<�XٕQP6@�4Μ�)�r��)�r��(J>�4� �@�������d�zAА000$O���������$ H�dɌI "I$000000e�	ɓ&L�2d��$ H��"��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	����"B�$�2dɓ&L� �e�	Y �e�@@"HI$��	�&L�0�"������������@�!�!�P�@l!0L
���9NS��9NS��9NS��9BPy�*�L"f��W,g��/$��a29�&rlDb���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�BK`� ���fJ���Z�?�$df�h�G�g)�r��)�r��)�r���X,Ca8㘘��"�T�C�@@ �"���������@�!D�&L``````�II !���A �&L�2dɓ&$H@�!D��"��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2dɓ&L��e�	�,`````````�I&L�2aD�������������Q(���H5��fY ��$�#�p �0�|�)�r��)�r��)�r���:)�c&��,	��28^Iy�ds0L�� ��e'��YI��@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���ʴFzVR+)?��X��3�@�V �2�* �f��9NS��9NS��9NP�|">d��<2�Tʑ�8G��/F�Y��2����������	L�2dɌI "I$000000H$d�A�L�2dɓ&L H�$O'������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	$H@�!D�	L�2dɓ&L�H2�	�,�2dɓ'�����������2d�  �)
F�؛8G������B�UF�!��3�,9NS��9NS��9NP�|
�|��``:eK�
�/32U�@F$�V
�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���ʴFzVR+)?�\pA �����&2`�4Μ�)�r��)�r��)���0������}>�
,�H�����������	L�2dɒ	X���$�$�A �&L�2dɓ&$O'�$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"B�$�2dɓ$�dɌ	X��������� �e�&L H��"�����������&L��@� d�#�p� l!0L
���3L�4 M�����}>�@�$T 3��9NS��9BPy�2A4lʨ�zn3Yl@�Ы@��3%PlDa�BK`���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����@Yc>���*؁=7��&2`0Y���t�9NS��9NS��9A�i�*�\������'�����������@�$ɓ$����������������,�H&L�2dɓ&$H@�!D��"������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H�$H@�!D�	$I2dɓ&H$d�A�H$c�A�L�0�"B������������L�1���t	�@�Ȇ]t�<�º!�0�3L�4%�)�r��f���$@(�2D|��)�r��)�� 8�!VE[$t*�<���Td��X+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��I�>�����.�B 3@�D���=�$A��4Μ�)�r��)�r��(�dp������"I�&000I$��	�'����������2dɓ&H$cɓ&L�2dɓ&$H@�?�	��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�2dɓ&L� �e�&L�2aD�	����������� H����Y��(
�#�`�b��4�3BPy�r��)�r��)�r��)�r��)�#L�	��V29�&rlDb���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����lDc#��g%䗐l tʗ��q�)�c&�σ��9NS��9NPX,eL��1
���/Dp�����G�6&�؃��H&L����������$ H�dɒ	X���$�$�@CY �L�2dɓ&L H��"B���	��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D����D�	$I2dɓ&L�2dɒ	Y �e�	Y �e�	Y2dɓ&$O������������"Ff�X�P(3&d̘���@�$�`�f��(<�9NS��9NS��9NS��9NS��9NS�� �3���A �W� �� ��*�YI��@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�BK`�<��g�:X�,2��6eTT��t�9NS��9BPy���y������$	@��U���`�$	��R*EH0�9D�Q'��������� H��"I�&e�	�H�I	Y�H$&L�2dɓ$ H��"B�� H����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	$H@�$ɓ&L�2d��,�2cY�H&L�@�!D�����������$```�k5���T������ ��4�*��r��)�r��)�r��)�r��)�r��)�r��(J>�U�pp�R�^Iy�ds0L�� ��e'�Q������O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O��@F#�V��z88#L��r��)�r��i�f��0L*
�8�> g)�r������$��yə3"�@��k5�&O�����������"I�&e�	�H�I	Y2dɓ&L�2dɄ	$O$ H�$O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"x@�!D�	L�2dɓ&L�2fY �000000000000000000L�2dɄ	����������� H����Y��P(�xg�? �~? `f��h<�3�)�r��)�r��)�r���X,��$!�0� �0Ca*
�8�9NS��9NS��9NPygFH&��a4dJ�$)S���� �� ��*�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O� ��*��A��̕Ay%��"���D���t�9NS��9NS��9NS��9NS�F��X,@(�?��(e�blM��!I  �"���������@�$ɓ2�����������������A �$�dɓ&L�2aD�	����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"B�$ H��"I�&L�2dəd�A�H$&L H��"�����������	e�	�D0�8�B���~6��~ �0��$�ʃ�r��)�r��)�r��(J>APga!�p0�G�3&d̟O������`�f���X,�9NS��9NS��9A�i��͐�	�����*^�g�:e�C ��*�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����lDc#��g&|3�,g�� ���H&���i�9NS��9NS��9NS��9NS��9NS����a0L  	���0g��T��a�rHL�?����������"x@�$ɓ$�@C�A�H$dɓ&L�@�!D�	$O����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"B�&L�2dɓ&L�3,�$I !���dɓ&L�2aD�����������$�2e�D�P(!���~6����<&	�`X,r��)�r��)�r��)��πX,!�0�q��3���2�2�
@@"I$_°a�r�T�����bł`�&��g)�r��)�r��)�r����S��L���M�	 JT��fJ�� ��$>L�+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�`� #Xφy�Xdp,G��g
p�ɀ�f��9NS��9NS��9NS��9NS��9NS��9NS����t��$�`��>�O�@��Y��L�?���������$H@�$ɓ2̲@������������2dɓ&L�2dɄ	$H@�< H�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$ H��"B�&L�2d̳,�H$d�A�000I$��	�&L�0�"�����������dɊ��|bU
�T2�P�2�Tʀ 	��r�FA`�Y�r��)�r��)�r��)���0�Î9�#��؛HR�  2d�� H����P(lM��>�O����f��!PT�A�9NS��9NS��9NS�d�h<���� �a��3>��Xd��X+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����2Ib�@g����K�e����T�HS��L6G)�r��)�r��)�r��)P| �S�2di{�P2F|�BS�*��r��)�r��)�r���X,Ca~?������g���)I /�����������&L� �e�I !���dɓ&L�2dɓ$�2aD�	��'�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������"B�$�2d�A�H$d�A�H$d�A�000000000I$��	�&L�0�"B������������L�1X�/�C���!��}2�Tʀ 	���0L��S��9NS��9NS��9NPM3���C  	��S*eO���6&�0�9D�Q'�����"EaX�
d̙�0�8��0L��S��9NS��9NS����tT#�08� ����Z���*�`� #����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�h�����2Ib�@g�� 
����� ��<�
p�ɀ�f��9NS��9NS��9NS��*�J|�0��6��M��2�2�=2B��
s`�&���T��9NS��9NS��9BPy�d��� @a @��3&dP(�f�d�����������$I2dɓ&000I$��	�,�2dɓ&L�@�!D�	$O��������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�< H�dɄ	L�2dɓ&L�H2�	$������� �e�&L H��"�����������&L�Q(�F�؛8G�2�T M���$��Py�r��)�r��)�r��(J>`�YW*�d M��?���2���0�9$&L��������2��P(Gdv��_��~?�03L�4%�)�r��)�r��)�T 1�	��>g�8dJ� � f��˦F2��!�BK`���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?����A	,U�`� #��� ���Yl@����N0,���:r��)�r��)�r��)�T 3�/�>l��,3@0 �32"��p �R��z4*�S
B �z��'͘� $g�č>
�P| �S��9NS��9NS�F��PT��������d�z�D�H H����������$I2dɓ&000000I$��$���� �e�&L�2dɓ$ H��"B�������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��"B�&L�2dɓ&L�2A �$�@D�H```�H2ɓ&$H@�?����������$I2d�$�:�� d�#�p� l%\���PT�(<�9NS��9NS��9NS�%� �X,��$3Fh��C(eblE!HR(�J$ɓ'�������$I2d���V(
d̙��xd�����g)�r��)�r��)�T 0,�
p�Ɂ�<�
�*؁/$��a ,��A��O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��V���J�FzVR+)?���͂��^fd��U�xS�� �$)�c&�hJ>S��9NS��9NS��9J��T 24�*�8F`�ffDA��T�d��	U*��G=9���F�z4sѣ�� J�T�h0'$|��9�p�ϛ!�*�P| �S��9NS��9NP�|�`��&	�sB!�
B��I$���'����������@�$ɓ$����I$000000000H$dɓ&L�2d���D������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"B�&L�2dɓ&L�2A �$�@D��I	Y2d��'�����������@�# �P(��G� @��!�0�3L�4F�Ӕ�9NS��9NS��9NP�|">d�0?���(e�T*�Pa�sY��000$O���������&L�$�!H��������~?a!�`�Y�r��)�r��)�r��(<�������X�,�f*�`� #����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�h�����VR6"1y���#�V�⬊� L�pp�����%�)�r��)�r��)�r��)P| ��ૌ�a�*�8_�|�@��h0' J�T��M�h�G=9���F�z4sѣ���h�G= �R��9/)��������d�&F���/�)�r��)�r��)�r��`�$G̐��TʙR8G�P(5��dɓ���������� H�dɒ	X������������ �e�	Y2dɓ&L�2dɄ	$H@�!D��������������������������������������������������������������������������������������������������������������������������������������������������������������������@�?�	$H@�$ɓ&L�2d̳,�L�1���I$I$��	�&L�0�"�����������	000�� ��G� `�� �0�3LД|�)�r��)�r��)�r���:f��h��G�����~6R*EH�P(��H������������AАd�z#�p�S*e@�<3L�4F�Ӕ�9NS��9NS��9@`�dlʨ�g���tʗ��K�6�����O�Z�=+)?�����O�e'��YI����VR+)?�h�����lDc#��g$t*�<���e������P����i�9NS��9NS��9NS��9J��F�\'���  ��2�2�	̈́����A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F����)���!_A�9�p�|r����)�r��)�r��)�f��h�g�����~6��"F�����������"I�&H$c�H```�H2ɓ&L�2dɓ&L H��"B��D�������������������������������������������������������������������������������������������������������������������������������������������������������������������	��$�2dɓ&L�2d̳,�H$c�H�I&L H��"�����������	I$���t$ ^�ə3&&&'��� �34�3NS��9NS��9NS��9NP�|">d�h�?���_��fLə
 �:?��������������	I �C�"�T�LLK,!�0���g)�r��)�r��)�r���:*���� �@�0 2!]6"1YI��@�g�Z�=+)?�h���@�g�e'���A�,^Iy�X�,2%\&3EB>	A���r��)�r��)�r��)�T 24�*�8M��  �zd�}����qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ�� J�Tʜ����@���~	��d��L�/a)���9NS��9NS��9A�i�	�`�q�1113&d̔
����'����������@�$ɓ&L���������������� �e�&L�2dɓ$ H��"B�'�����������������������������������������������������������������������������������������������������������������������������������������������������������������"x@�!D�	$I2dɓ&L�2dɌd�A2dɓ&$O�����������ɓ&
�P�E�_��~?�("��3�`�Y�r��)�r��)�r��(,3L�4�QX�`0�fLə
�Y��$�����������������D�&L�k5� ^�P�G��� �34�3BPy�r��)�r��)�r��(l��UX#%��2��*�Xd��X+)?���͂��e�F|3��Ҧ#�U	�L�N0�|�)�r��)�r��)�r��A�	O�p�b���zd�}����qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�l%T��,�A6fdf
���t%>��/�)�r��)�r��)��ρPT�����8G�I�����H���������� H�dɓ&L`````````�I&L�2dɓ&L�@�!D�	���D�������������������������������������������������������������������������������������������������������������������������������������������������������������$O$ H��"B�$ H��"I�&e�d�A �$�������������dɄ	$O������������&L�@�P111��<�3L�X,T 3��9NS��9NS��9BPy�f��h��q� `�d̙�@�Pk5��$�2d�������������������"I�&Q(�CC�"�T��3� �L��X,�9NS��9NS��9NP,�
�|FFh&�?�$t*�<��U�|3��%*b�#�U�y��1��͐<�3�)�r��)�r��)�r��A�>
��	@1�,)̀g�HWњ)�P8
 J�T��M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���%T�eNFK�e e�\�6��&���T��9NS��9NS��	A���*�U�ɑ��+��_��Gdv���$�&L�����������D�&L�H2�	$�$�&L�2dɓ&L�0�"B�$ H�$O������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	$I2dɓ&L�2A �&L� �e�	Y �e�	X@�!D�����������$�2fY �e�	D�	�@�P�C(Car��)�r��)�r��)��πX,�0�@�"te� d�(
(�J$ɓ���������������������"I$�(
6&�،��2������Tq�r��)�r��)�r���4Ό�M�2�*�<��&i�*����xJ>S��9NS��9NS��9J��T 1�6B����&zd�}�S���%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��X&�l���  '��J|�)�r��)�r��)�r��`�$G̐��TʙS"teҁ@�001����������$�2dɓ$�@D�H�I	Y �e�&L�2dɓ$ H������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�$H@�!D�	$I2dɓ&e�d�A �$�dɓ&L H�������������$�t$
��T��#�p��8Gdv���)J%T*�P����(<�9NS��9NS��9NPX,Uʹq� G�6&�؊B��I ��'����������������������2d�f�X�P(2!�F] `� l&H�� �|�)�r��)�r��)�r��)�r��)�r��)�r��)�T�J��a�*�ٙ�) #/*r2^P��L�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѠ	U*����f
�S� �3�% ς���)�r��)�r��)�f��h�fTʙQT*�QD�Q�����������$I2dɓ&000000000000000H$dɓ&L�2d��$ H�$H@�?�������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�	$H@�$ɓ2̲A2d��,```````````````�2dɓ$ H�����������$```�k5�
 B!�����?���x�P
 @(&F20���0g����eL��2D|��)�r��)�r��`�!�0 �	�2�T�}>�blE!HR(�J!D�������������������������J%HR�P�E�_��	@��#�H�> g)�r��)�r��)�r��)�r��)�r��)P| �|�!8M��  p��x�����*�S7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aҧ#%��/�>3@	��:� �P| �S��9NS��9NS�Tq��~6&�ؓ&O�����������$�2d�A�000000I$��	�,�2dɓ&L�2d��&L�@�?�����������������������������������������������������������������������������������������������������������������������������������������������������$ H�$H@�!D�	L�2dɓ&L�2d�A�000000000000H$dɓ&L�@�?������������&L���k1Gdv�(e����3Fh�f��(<�9NS�%� �X,��$d���	A���r��)�r���� �3���}>�H��R�"HL�?��������������������������ɓAАfLə @a��t�9NS��9NS��9NS��9NS��9NS��*���W3M��f
�f�p��L�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U1�	�	 �)̀3�e�|�'�P_�S��9NS��9NS$G̐�C(V/���@�!D�	����������@�!D�&L`````````�I	Y2dɓ&L�0�"B�$ H��"x@�?��������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"B�$�2dɓ&L�2d��,``````�H2��,�L�2d������������$�$
%��``lM��>�O������$G̐,9NS��9NS��9NS��9NS��9L�4� @��6&��k5�d�G��������������������������L�2I$k5�́�/C(e�<�Py�r��)�r��)�r��)�r��)�r��)�	@08_�|f�p��Lsѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�@�(D/@p���  ɑ���*��r��)�r��(<�2�Tʔ
���I$+
��(
�!H0�8�``+�����2d����������@�$ɓ&L�$�$�@D�H`````````�2dɓ&L�2d��'��������������������������������������������������������������������������������������������������������������������������������������������������� H��"B�$�2dɓ&L� �e�	Y �e�I !������,�$&L H��"���������� H�dɒI  P(lM��>�O������U�Ȩ*��9NS��9NS��9NS��9NS��9NPX,8�O��@�PQ(�B�������������������������� H�,�H5��a&`jdC.�� ���da]�C�`���9NS��9NS��9NS��9NS��9NS��*���*�i�D/A@�(�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���	U/���zd�}6c$ ��8r��)�r��( �	��}*EH��8G���������~?���2fL�@�P$��Dɓ'��������� H��"I�&H$c�H�I&L�2aD�	$H@�!D�	�������������������������������������������������������������������������������������������������������������������������������������������������"B��D�	L�2dɓ&L�2dɓ$����I$000000e�d�dɄ	$O������������"I$��)
F�؛���@��Caf��i�r��)�r��)�r��)�r��)�r��)�r��)�f������2�Q�6&�BA2d������������������������	H$f�Y�P(�2fLLLO����fH�� �|�)�r��)�r��)�r��)�r��)�r��)�r�A~���� #8��L���4�%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M����D/@g���8r��)�r��)�f����x@(�	�`��3L�X,��`�Y�#�H�����2�P�6&�؂�@�����"���������@�$ɓ$����I$I$��	�,�2�ɓ&L�@�!D�	$H@�?�����������������������������������������������������������������������������������������������������������������������������������������������"$ H��"I�&e�d�A �$�dɄ	$O�����������dɒI !B02@��8G �3�bń0���X,�9NS��9NS��9NS����tS���A #>e$d��F�Ӕ�9NS��9NS����t&	�`H��������#������������������������e�	�Y��P("�T��g�`��� ̑2G)�r��)�r��)�r��)P| ͑�0YU�Qx8 � �r��)�r��)�r��)�� �N�ј*�8_�|D/A@�(�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���hUJ�T�d��R F^�O��PHϑ�P| �S��9NS��9NS��9NS��9NS��r�FK,bbbT��R(
�|_&O����������	L�2dəfY ```�II !������,�$&L H��"B�'�	�����������������������������������������������������������������������������������������������������������������������������������������������$ H��"I�&L�2A �$�dɓ&L H������������ɓ$�@@�:�A�3&d��ıb�C`X,�σ��9NS��9NS��9NPygE8�>
��#G	���� W���2f@�@ϊq�|�)�r��)�r��(J>�2C�9����B�R�"�D�$O�������������������D�	Y��k1*�P�>�O������$G̐,9NS��9NS��9NS��*��2fh,�����"��9����E���l��� ��)�3�fT 3��9NS��9NS��9J��	@1�,)̀^`�Fh0'6�_�qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�@�(e�a��&�̀�b3�e�|�%A�*��r��)�r��)�r��)�r��)�r��)��σ4�3Fh�2�Tʑ�8G��/@�P(``` H����������$I2dɓ&000I$���,�L�2dɄ	$H@�!D�	�������������������������������������������������������������������������������������������������������������������������������������������� H�$H@�$ɓ2̲A �e�I !���A �&L�@�?����������ɓ&000k5���AR*EH��ıb��4�3A`�Y�r��)�r��)�r��(<�3��d�1~	J��ɟ�/�~^#� g�����ʘ���/b���E`���+��S8@ϊq�|��:r��)�r��)�r���:f��h��FTʙR�T��a�rHL�?�����������������D�&L�
B��lM��>�O������$G̐,9NS��9NS��9NS��*��$h&��8��� ��=	!T�٘�&@�B��`N$��j6B/)�F@��i�ȑ�� �r��)�r��)�r��)P| �S�	��:3@0g�HWі	�Bl%T�����z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���	U/�����0�6 ���% ς����9NS��9NS��9NS����dd��dd���2NS��9NS��9NS����e\���]21��LLA�x)
B�$&L����������$�2dɓ$�@D�H```�H2̳,�L�2dɄ	$H@�!D�	�������������������������������������������������������������������������������������������������������������������������������������������@�< H��"I�&H$c�H�I&L H������������D�	Y��k(
H�#H�02D|��`���9NS��9NS��9NS�F��M3��*s�&��x���&��&}�iE0^�#@��Q�(�h��(��>)�X2��ʹ�r�e$d)�I�#L��r��)�r��)��σ$G̐�g����}>������'���������������$I2d�@�Q�6&��}>�S*e@�J�W#"��3�Py�r��)�r��)�r��)P| πx�#A4�LU�0� �$�R*b��:P2a���I`N$�2"PȉC",	ĕ@�F �@�^��	1�!>l��UDM��2����)�r��)�r��)P| ς�� �P�3�0�6����9/)��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSM�M*r2^S) #/��'��?�24����8T 2����)�r��)�r��)�T 3dd�М�p��R�U�g*�Xq�F��1l���r��)�r��)�r��(,2D|�њ?�ϧ��2��k5�&L H����������$I2dɓ&000000I$��	�,�H2ɓ&L�0�"B�������������������������������������������������������������������������������������������������������������������������������������������� H��"I�&L�2A �$�@D�A�L�?����������$�2f�Y��P("�T������~?�xd�����g)�r��)�r��)�r��(<�3�1~	J��ɟ�/�~^L�O�h���>`hB4
!��F�D#@��Q�(�h�G��5S&�(�̫��F�Nzd�b���)�r��)�r��)�*
�8 �3���2�P�6&�؃��H&L��������������񁁀P(d�z#�p� @�b���	���9NS��9NS��9NS��> dh&��8�B��� M��4�&�E�	(W�|X�%��2"PȉC"%��2"PȉC"%��2"��HIB��AxB<��8�*b�#A4*��r��)�r��)�r��A�������3�$+���	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M
B �z��'�`�p�ϛ!�*��r��)�r��)�r��)�l���6bf���V�f��g�	��rV_�9+/�g�@�OW713��Pϊ�1�r��)�r��)�r��(�*�
D$	E�_��@�3���H H����������$H@�$ɓ$�A �$�dɓ&L H��"B��D�����������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2d�H�II !���d�����������ɓ&k5���!�P�G�����$G̐<�3�)�r��)�r��)�r��(<�3�1~	J��ɟ�/� g�8fPǀ4/.L��:�`��<���L�04
`h��(�hB4
`h��)��Q�(�h���/gɴD̠!��#��BpL_�PygNS��9NS��9NS�F�ҮU��$	E�_��*�P���A#������������D���H	0�S2fLɉ��$	@�PT�)�r��)�r��)�r��(J>�Mq��6e���0��J�'*�0
%�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"�����F �<�(�7YU6FL�9NS��9NS��9NS��>
����tٌ� �O�HyS���"�9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�AРp2�0�L��
�)̀)�`l	@3�/�)�r��)�r��)�r��)�2fh,و�z+�W71	�" L�(3�����e��}.?K��������C(�#��^�&GeT� �3���8/f�ə�)�r��)�r��)�r���:d��� @a @�#�p���� �2��������� H��"I�&H$cɓ&L�2d��$ H�����������������������������������������������������������������������������������������������������������������������������������������@�!D�	L�2A �$�@D��	���������$I2d�%�a�r;#�D>�O�TʙP<̑2@�X,�9NS��9NS��9NS����t&/�)���$� �#�C2��<�xrg�f��S���)�<�৒<��)��S@��L�04
!��04
`hB4
`hB4
`h���/b��=>�¨��,��)�r��)�r��(J>�4� @a/��/�B!�
B��Q(�B�����������D��f��@�T��R/��/����@(�A�#L��r��)�r��)�r��)P| ��MeTD�7�2����� NU�`Kq%�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'X�*�0
%N "�
U� Bx�N2��h&���<d��)�r��)�r��)�T 0J�pX
s`>C4�%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�l%T��4�Hx/�>l�H 2di{	O�p�> g)�r��)�r��)�r���<d��8f�^ Fa������	���!��e��}.?K��������}.?K��������}.3�3	�����@ !�2 p��Q�+�	�aP| �S��9NS��9NS��> `�X,�Q~?�P�DvG`�)
B�$&L����������$�2d�A�000000I$��	�,�2aD�	$O���������������������������������������������������������������������������������������������������������������������������������������� H�dəfY ```�J%����"��������L�2H)
B��6&��}>����<̑2@�X,�> g)�r��)�r��)�r���4Ίq�|I�T �3����eɟa�GQL�@��O$x)�04
`h��)��S@��L�04
`hB4
`h��)��S@��L�<�৒<�G���S�eɟa�)�X3� 
��r� ���$���t�9NS��9NS��*��f��4f�S*eLə3%�@�Q(�&O���������2���D�bU
�T_��_���� �34�3A`�Y�r��)�r��)�r��(J>��0x8 ���"F@����� NP����B0J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8������F �<�(�74A�dg��9NS��9NS��9NR�����8d���l�H M��`�d!@�(�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSM�M
B �zM�����x	O�p�> g)�r��)�r��)�r��A�#Bp��1d��R�9{ ��b��Q�L�2��~>������q��\~>������q��\~>������q��\~>��e��C(�#��^�&Gb	���_�E�1|�I�r��)�r��)�r���X,��$��y�eїJ���k&L�@�?���������D�	L�1���I$000H$dɓ&L�@�?����������������������������������������������������������������������������������������������������������������������������������������	$I2d��,```�Q(�@@"d���������@�$ɓ$�@@�P(؛b}>�L��2�l"CaPT�(<�9NS��9NS��9NS����tS���A #>	3�0�0U�QL��(��>j2�04
`h�G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�S@��<���/c.L����(�̫��/�`b�d�)�r��)�r��)��σ4�3@0?������P(��L�?������	$ID�Q�!HU
�Tg�? �?�њ�0,9NS��9NS��9NS��*�� �pA3M�D&�r��x��P@�B��`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%P2�:P2�1�LA6O��� �Qdg��9NS��9NS��9NR���A~�����W3M�R F^T�d�����z4sѣ���h�G=9���F�z4sѣ���i��)�	U*����L����8Xg͐�|��> g)�r��)�r��)�r���ə��f K���\��e�� L�(3�����e��}.?K��������}.?K��������}.?K��������}.?K��������}.?K�#>�&bFa3����d^DU���eBp8^͑�3J��r��)�r��)�r��(<�3L�4�Q	@��C(؛b
�����������$�2c�H```�H2ɓ&$H@�!D��������������������������������������������������������������������������������������������������������������������������������������� H�L�2dɒI "�D�I ��/�������$H���(
6&�ؑ�8G 8�a!��4�9NS��9NS��9NS��9A�i��͑������@0�0U�PE� ���E0^��H�S�
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��H�S�
`h�eL|�DE\�Us96c������)�r��)�r��)�r���� �@����2�Q�6&�BA2d�����D�J%HR����}>����6�U��,9NS��9NS��9NS��9O�x���	�n2!0�L���I
�T�R/F��T�`�'J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DX�*�0
&�E�# A�a��G3M�D��p%�)�r��)�r��)�r��g͐�3�e�`���
�3A�3 J�T�=9���F�z4sѣ���h�@�U1�	�	 aNl�d��L�/a)���9NS��9NS��9NS��> c>*�pUBJ�1 ��2"����g%e�3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������p$g�D�C(�&�`4��<*�Xr�z+�,و����)�r��)�r��)���`�&q��3���2�P((�J$ɓ���������@�$ɓ$�@C�A�L�2dɄ	����������������������������������������������������������������������������������������������������������������������������������������"B�&L����$�/��X�	������$I$��F@��8G቉�bŀ("��3���r��)�r��)�r��)�r�q�|I�T �3���"�B�#��ف�S�
y#�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�S�
y#�M@�T�ɴD̠!��#�#
�\���4Μ�)�r��)�r��(<�3�\���H��������!HR��ɓ&I �!HR6&�ؑ�8G 8�r�FA`�Y�r��)�r��)�r��)�|�H<FqS`	�	�B|�x7<J�d#�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%�8�s��x�Q�,_�YU6Fpl�S��9NS��9NS��9O���24��1�  �~	�) #/*r2^SqSG=n �hUJ�T�d��R F^�O��PpWF|�%A�9NS��9NS��9NS��*��`N��#�&r*�{ ����P3����F}�$O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����1�0��Y���������ʄ�p���8f�)�r��)�r��)�T 34�3@0?������؛b!	���������&L```�II "A �&L�@�!D�	�������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000I �%����@�?������$�@@�:�A�3&d����!!�0�*�ygNS��9NS��9NS��9A�i��$�@ώ"���M��� W����"�p"GQL�@��<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!��H�R:�`����Dx@�@� �p ����t�9NS��9NS��9BPy�d���q�LLA�x)
B�$&L�2d�  (
	0�S2fL�x21��t��r2��Py�r��)�r��)�r��)P| πx�#A4	�Rٖ/� 2��g�a"�@�Fq$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$��(��R�zB��� 	�R��p�����9NS��9NS��9J��3��A�2����Iє�����S� g ���J��r��)�r��)�r��)��σdd��Y�%��W�nb2�Q��&�Y�#>�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\f!�f9+/����OW713��P,و�2NS��9NS��9NS����fH��!���ĩ"�P(
%�2d���������	Y$�$�@C�A�L�0�"���������������������������������������������������������������������������������������������������������������������������������������"I�&H$d�H�/�b�D�L�?����@�$ɓ5��e�@�"�bbb	@� ��3L�X,r��)�r��)�r��)�#L�'�L_�R�=2g��� W����"�p"j2�04
`h��)�<���L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�F�D#@��S@��F\�����S? �AL��H�S���F�Ӕ�9NS��9NS�F��4�3@02�Tʙ�2fL��/F@���T�����bń0� �3��x�9NS��9NS��9NS��>�$��pUDL�q��Q�l#<��(��Kq$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�'nx<�� �\e���q���	�2fiP| �S��9NS��9NS��> a)�24���aPU 0�>
��T 3��9NS��9NS��9NS�2F|T	�p�  �{2��dE\�L�f�����C(�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��e��C(�&rV_�<�ϑ�EZ�`_�Y�&�ə�A�9NS��9NS��9NPX,f��h�g����}>� ^��t$I  �"������$�H2�%�$�&L�@�!D�	�������������������������������������������������������������������������������������������������������������������������������������@�!D�	L�1���I$+
��$'�����"Mf�Y��"��$	@�">d�`�Y�r��)�r��)�r��(<�3��4΄��%*s�&��x���&�P!�1��S@��Q�(�h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��H�S�
`heɟa�xB�*�
��ɳ# 8�$���t�9NS��9NS��9EAPg P
 Gp6
D	�#�H6G)�r��)�r��)�r�����dd��YU6e���0��J�'	(W�|U!%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��IB��@*��� ��)�2fi�r��)�r��)�r��)P| ʃ�r��)�r��)�r��)P| ʃ�F�����3����dE\/3�s��2��	� �?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3	��Q�M��(��add3���%>Ô�9NS��9NS��9J���ʹW#&F20�����"�T�C�J%d��������dɒI "HI$���,�2aD��������������������������������������������������������������������������������������������������������������������������������������&L�2d�	  �+ĒH H�����f�Y#�p�b�0L�`���9NS��9NS��9NS�F�И��Nzd���? �&g��4/.L��:�`��H�S�
!��04
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)�<���F\����4/�@���F�Nzd�b����:r��)�r��)�r��(<�9NS��9NS��9NS��9NSdd��YU3M�D������@(��"��I(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���J������2��x�����q�#A49NS��9NS��9NS��9NS��9NS��9NS�2Af�@��0/�U*�3����3���J��f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3�!��	��xW�`_�Y�'�P_�S��9NS��9NS����t��$��y�2�T�}>� ^��t$&L H������ H�����D�I �$�2d��'�������������������������������������������������������������������������������������������������������������������������������������$H@�$ɓ(�J&�Y�``` H����L�3blM�błPy�r��)�r��)�r��)�#L�L_�R0�����@�����eɟa�`hB4
y#�O$x(�h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x(�h���/gɟq��0�D'
q�|�)�r��)�r��)�r��)�r��)�r���34&i�Ȅ�=2�J�@J��E���y*����DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DX��e!�l�����9NS��9NS��9NS��9NS��9NS���1�*"�D ��Pg%e�3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFa3����d"�DF@<�U	(g�@��9NS��9NS��9NS��a!� H/��/�T��a�rH$O�����dɔJ%���$�2dɓ&$H@�?������������������������������������������������������������������������������������������������������������������������������������ H��"B�&L�$�(�J&�Y�``c����HG� �@��)�r��)�r��)�#L�L_�PH)��@ૐ*��4/.L��@��D#@��L�F�D#@��Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�S�
`h�eL)�X �33�)�r��)�r��)�r��)�r��)�r� �*� '��I
�T�R/@t�d*�0
$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$��(��$`3��? dg��9NS��9NS��9NS��9NS��9NS�g
�"�Dg%e�3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFa3�3�!��	��U*�3�"���f M��3NS��9NS��9NS��	A���f��x� @��8(
f�Y2d�����ɓ$��E�|+@@!���dɄ	$O�������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$�|_
ƳY��I	����  ��}	�`��9NS��9NS��9NPygG	��e�\��S�B4
!��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��(�hB4
`h��(�hB4
!��H�S�
y#�L��S��eL|�DH��韁 W��*
q�|�)�r��)�r��)�r��)�r��)�l��ـ� T�R/A%
�/�q$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DX�3�L�~�a�1*@���# ns4�dH�M
��r��)�r��)�r��)�r��)�r��)�3�L3���!<d@	��rV_�1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��e��J��F&G3 �����0/�Nٲ2fiP| �S��9NS��9NS�%� �X,Ca	@��C(P(����$���k$��Cɓ&L�������������������������������������������������������������������������������������������������������������������������������������'�	L�2A �$�@B��_�f�I$����D�Q>�O�\�����9NS��9NS��9A�i�@ρ���1��W��#��؄h�G��F�D#@��L�04
`hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
!��04
!��F�D#@��L����|	�"< zg�@������L�L_�QN2O���9NS��9NS��9NS��9NS��9NS�2FqS` 2��@E%
�/�q$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DX�,	ĕa�a"� �d��f���,���#86g�<d��)�r��)�r��)�r��)�r��)�r��)�l���6b��6L�U�<�ϓ9+/���Q�O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��2��g%e�73�^�&GeT� �_�E#Bp�9NS��9NS��9NS����e\���*eL��P(&L����$```�k5�J%I$H$aD�	�������������������������������������������������������������������������������������������������������������������������������������@�$ɓ$�H+
���k$�@AD����H}>�J�W#')�r��)�r��)�r���4΄��%*s�&�rl�\�U>M�$u�{04
y#�L�04
`hB4
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L���F�D#@��Q�(�hB4
GQL�E
�D`E�	�� W���M��!8A #>)�I�#L��r��)�r��)�r��)�r��)�r��)�r���ə���"l��D`3�(q$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJT�`��y# A�`���?  �e!A���|�I�r��)�r��)�r��(<�3�1~	D3�1~	A�i�9NS��9NS��9NS����Y�%��W�nb2�Q��&�Y��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����1�0��Y����W����3NS��9NS��9NS��9NP
D	��}(�J?����J%�D�I$���,�2aD�������������������������������������������������������������������������������������������������������������������������������������$I2d�	  �+ƳY��I���I ����W*�d�9NS��9NS��9NS��9NQN2O�0������"�*�4/�C*c@��<�G����F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x)�<���SP!�0"�p"�"�ϸ # ng&̪h� ���$�9NS��9NS��9NS��9A�i�2D|� `��x����)�r��)�r��(J>�M�q�# nr0�C @�F	C"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��B0@�B�@*�	�ze�7x8 � �r��)�r��)�r��)�#L�'����$� �#�? ��@�$�����8�>S��9NS��9NS��9M��3Bp8^�a�������|��Y��2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\f!�f�2�,l�	�r��)�r��)�r��)�f��i�t$���000Q(�J%�$�$�dɄ	��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�H2�$�|_
ƳY��I	����  ��}�C�)�r��)�r��)�r��)�r���d�RF@g���p FE2+ �.L��@��Q�)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��Q�(�h��)��Q�(�h��(�h�G��H�Q�)�ʘW��Ȭ�D^e\0��������'�<�3�)�r��)�r��)�r���X,��$�`$	F&&&d̙��T����}?���x��i�T 3��9NS��9NS��> f���N2��0�L���4#�bT�9V�Q,	Ē�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���BJ�_�R�`3�WplfX����"|�I�r��)�r��)�r��)�)�I� ��20��rl̢/2�)�Xrg�f����\�����S? ��/�Nzd�b����:r��)�r��)�r��)P| �f�@���_ʩV���L����(�e��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3	����EZ�P&9NS��9NS��9NS��9EAPgS*eA@�W�����Y��Q(�I "A �&L�@�?������������������������������������������������������������������������������������������������������������������������������������D��"I�&H$d�H�/�cY��I$�����$�@Dp��
D	�r��)�r������2NS��9NS��9NS�F�� ��$���)�Xrg�f��S��G��H�Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��D#@��Q�)��Q�)�<���S@�u�{rg�f� м�0a�	3�)# 1N2O�ygNS��9NS��9NS��9BPy�f��h����F�0�fLə
�Y�```�$	  a�s2fLɕ2�T��4�3BPy�r��)�r��)�r������Q�~  �D�J�'*�0
%�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'U!7<Fi>D`���?  YU6Fplʃ�r��)�r��)�r��)�� ���`g��� W�\@�(W$u�{#��ف�S@��L��S�B�L�@�#�#
��N2O���9NS��9NS��9J��F�����+�b!<d@	��rV_�1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\f!�f9+/����F+�b8/eA�9NS��9NS��9NS��9EAPgS*eA@�W�����Y��k5�I "A �&L�@�!D�	������������������������������������������������������������������������������������������������������������������������������������$H@�&Y�H$�@E�|+�f�I$$O���$�@Fd̙�
D	�r��)�|�HN2��i�Ȍ�*�x8 � �r��)�r��)�r���4Έ gʠg�@�"���_|���/f�D#@��<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�(�hB4
y#�D#@�u�{5S м&g� g�8	3�)# 0����d�)�r��)�r��)�r���4΂�`��&	�rˣ.��I��:��HL�0�"�ɓ$��B���B���� M���$�σ��9NS��9NS��> f�ə���"l��A6O��1�L$�_��`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%P2���~�N "�
U� Bx��*b�#A46FL�9NS��9NS��9NS����tS����H�
g g�8  ��� м�3�3H�)��!04
`h��)��S@��O$x)��R:�`����@�. L���I�q�|��:r��)�r��)�r��)�2fh,و$^ ت�`����WBHy3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFaѐL��쪕`̑x`Y�&�ə�)�r��)�r��)�r��)�r��i�eL���_��� H�,�$
±|k5��$� �e�&L H��������������������������������������������������������������������������������������������������������������������������������������@�&Y�H/��X�k5�I /����ə3 ���9NR���ʨ� 2��g���x�����q�#A4*��r��)�r��)�r���:Ȗd`!P0�#� g���E0^�$x)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
!��5S(W"	���AL��L�L_�QN2O���9NS��9NS��9NS�%�0L8�#�p�blD#�D�L�?����#blM����l H�`�&	A���r��)�r��)�r� �4�d@��F �<�2���'J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8��3 �F%H��4#�d��f���,���#86eA�9NS��9NS��9NS����t��"4q�f
��)�Xrg�f��S�B4
y#�O$x)�04
`h��)��S@��L�H�S�
!04
2�ϰ�<�xrT0�20�Ȗ#L��r��)�r��)�r��A��P&3��Q L�2�Q����L�e��C(�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��Q�L䬿�	��!<dB�F 3�x�1|�I�r��)�r��)�r��)�r��)�f��i�2�T
���000+
���k$�@Cɓ$ H�������������������������������������������������������������������������������������������������������������������������������������$H@�&Y�H(�J%�|+I  �"���$�3&d̀`r��)�T 34�dH�g�s��C 8����2��i�Ȃʨ��')�r��)�r��)�#L�L_�Q�Bpa�fP�ɴD�eL`h�G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��H�S�
!5S9�D����x��َ"���#@`�dr��)�r��)�r��)�r��`��&	��L��2������C�J%d��������2`�:��6#(e����@(���g)�r��)�r��)�T 24A�4�dH����x EP�P2���I(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$��(�!��xM��̱�q��6Fplʃ�r��)�r��)�r��)�#L�W2DiS��073�fg�@�< z�\��S���)��S@��L�04
`h��)��S@��L�04
`h��(�hB4
`h�eL�\�&g� g�8	3�0��N2O���9NS��9NS��9NSdd�М��F�/"*�yy�"�Cɘ�Q�O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����1�0���L���`�a�l�	�2fi�r��)�r��)�r��)�'�<d���9NS��A�eL���_����	Y��k5��d�```�2aD�������������������������������������������������������������������������������������������������������������������������������������$H@�&Y�H(�J&�Y��I	����$��3&d �3��9NR���2��# A���s����y EP�bT�9��fX����"l���r��)�r��)�r���4Ίq�|9� �3��6������H�S�
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x)�<���M@�T��mXqg� �73�f8�N*�H��$�9NS��9NS��9NS��9A`�XL�4f����?�� �C<1Q(�I�'��������ɓ(�J"�@���8eL���4�3L�ygNS��9NS��9NS����	�R&�r0�C @E�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��(
��E��BHU �qSa	��P| �S��9NS��9NS��9A�i�	��JF p	3� 3�L�O�h��ʘ��)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��Q�)��Q�&}�h�E`�"�*����S��0����4Μ�)�r��)�r��)�T 0Y�&H��U*�3����s��2��f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��2��g%e�7 �	�"*��#8W�dd�Ӕ�9NS��9NS��9NR���#86a8�B�2���� ��)P| �S��9L�4�2�Tʂ�@������,V��Y��I$���A �2dɓ��������������������������������������������������������������������������������������������������������������������������������������&L�2c�D�k5�I /����
�R*@��)�r���70���y�e!���nx<�� � �J�'# A�`���,_�YU6Fpl�Py�r��)�r��)�r���:)�I�F p�rl������eL`h��)��S@��L�04
`h��)��S@��L�04
`h��)�04
y#�O$x)��SP!�0��>)�XrT0�20�Ȗ)�I�r��)�r��)�r��)�r��`�$G̐�g���������R*E�@�Q(�d�@@�?���������ɓ$��A�!�ə3$��<��$�σ��9NS��9NS��6Fpl�eTDf� *�#�	�J�_�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'X�*�0
$bT�9xB<F@��i�ȃ���������)�r��)�r��)�#L�'�� F|��B�a�*�
���˓>�4���/f�L�H�Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
!��F�D#@��C*`E
�D@A3=>�¨��N2O���9NS��9NS��9J��l������+�b!<d@	��rV_�1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��Q�L�2��nf9@��L�ʩV���6�1|�IP| �S��9NS��9NS��> g�<d����7�g�Q��g�a"�!����6	���r��(�*�*eL�(
����```V��Y��I$��	�&$O'������������������������������������������������������������������������������������������������������������������������������������ H��"L�,�000Q(�Mf�Y$�'����
�T*�09NS��*��n2$`3����nx<��&�ɹ��nx<�� � �J�'�p�M��0� q��6FL�*��r��)�r��)�r�q�|I��/�Q�W<�x5S04
y#�L�04
`h��)��S@��L�04
`h��)��S@�u�{rg�f� м
��f@�3�d� �4Μ�)�r��)�r��)�r��f�Tp���#�T���P(5��cD�����������$�I
B��@�3�6$G̐<�3�)�r��)�r��)��h,���2���Q{3$�J�_�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'U�`@T2��fX����"l��ل����9NS��9NS��9NS�F�И��Nzd���>� ��dVE|	�":�`��F�L�H�S�
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�F�D#@��Q�)�<���R:�`����B��S? ��/�RF@b�d� �4Μ�)�r��)�r��)�|�l�	�/ l �ȫ@yy�"�Cɘ�Q�O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������C(�&rV_�129��dE\/fTg
�3�L|�I�r��)�r��)�r��A�6Fpl�q���� g�$*�{3$��@�U!,	ĕ@�F )V�<NS��9L�4�2�Tʂ�@������,�k5��f�I$e�d�dɄ	$O���������������������������������������������������������������������������������������������������������������������������������������2dɓ(�J&�Y��	�����x�`�r��)�f��������s����y7<M��s����y7<M��s��J�'*b��=	!T�O�LU�h&��A�9NS��9NS��9NQN2O�)# 0H)��xS"�
2�ϰ�04
y#�D#@��L�04
`h��(�hB4
y#�D#@�u�{rg�f� м
��fAL�� �,L�g��i�9NS��9NS��9NS����t�a!� H1113&d̊�t	�H H����������������F�؛?�� �$	�0L��S��9NS��9NS����x8 ���"U�\ f������r)���PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC",	ě�%LU"� �'�a� �)
�2NS��9NS��9NS��9NP���`g��� W�3���"j2�#����<�৒<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)�<�৒<��(˓>�4���̠!��#��Bp� F|F�Ӕ�9NS��9NS��9J����pUBJ*��"!<d@	��rV_�1�0������q��\~>������q��\~>������q��\~>������q��\~>��e��J��nf9@e��*�Xs$^ �l�	�2fi�r��)�r��)�r��)� ��"f���Wpl0��A��XfD�'J(dD���@)V�<NS��9EAPgS*eA@�W�����Y��k5�I #,�H&L�@�?�������������������������������������������������������������������������������������������������������������������������������������	$I2d�
%���k$��AD���񁁀B!�њr��)�r���""m#s����y7<M��s����y7<M��s����y�e!���l �^R�*�z3ВH ���T�XF�h8T 3��9NS��9NS����tA #>	3�? �,���'���)��y#�O$x)��S@��<�G��F�L�����h�!�@C�@��r�T�L&/�(<�3�)�r��)�r��)�r��(,�C,X�<�8G��6"�`I$������������������&L�:��blM��C(�?�P
 A`�Y�r��)�r��)�r����pg1V�79� ���
�d#���DJ(dD���DJ(dD��@�F �@�T�(/ hG�a��G3M�D'�<d��)�r��)�r��)�r���d�RF@`�S8 �3\�U<�x�'���)��y#�O$x)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�S�
y#�H�)��+�O�� 3� 3�����X�'��r��)�r��)�r��)�2fhN��#���p<�ϓ9+/���Q�O�������}.?K��������}.?K��������}.?K��2��g%e����/"*��{2�8W�4'Ô�9NS��9NS��9NR������)
 Bx�����E��`��e!`N$�2"PȉC"%��2"Pȋq&zB����9NS��3L�*eL�(
����```�k5��f�I$e�	ɓ&L��������������������������������������������������������������������������������������������������������������������������������������D�	L�1����D�k5��%�@�?����$P�C4f��)�r��i�ȗ�4#�� ��y7<M��s����y7<M��s����y7<M��s����y6B/)S����	�ze�7x8 � �r��)�r��)�r���4΄��%������ 3�E
�D���/f�D#@�u�{5S&�< zg�@������L�L_�PygNS��9NS��9NS��9NQPT�C`6*eL���}6&�؂�@�I$L�?�����������������ɓ(�J"�@���8?���<2D|���:r��)�r��)�r�����N2��0�L���4#�bT�9V�Q,	Ē�DJ(dE�8���~��E�# A� ��l��UDM��3NS��9NS��9NS��9J��)�I� ��D'���3? �
dVE|	�":�`��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)�04
`heɟa�xB�ey�p73�fT�L&/�(<�3�)�r��)�r��)�r����l�	�/ lUJ��4��<7 �3�����e��}.?K��������}.?K��2��g%e�7 ����W712E��f�@���9NS��9NS��9NR���#86`��"f���p3�� ��E�*�0
%�8�PȉC"%��2"PȉC"%��2"��IxB<��9NQPT�TʙPP(������b��k5�I !���dɄ	��������������������������������������������������������������������������������������������������������������������������������������$�2dɓ(�J&�Y��Q(�	���������9NS��7��x��y7<M��s����y7<M��s����y7<M��s����y7<M��s���A��N "�h!�79�n2 �pA6FL�9NS��9NS��9NPygBb��"��#����6��&}�A\@��x�9~*s�&��F��ygNS��9NS��9NS��*�,	�`������2�P�6&�؈F�D�2aD�������������������dɒI  ��d̙�*eL���H�� ygNS��9NS��9NR���#&f�ʨ��?  
U�F%H��2����j7<J��E�A6O��� 	�R����͑�r��)�r��)�r��(<�3�1~	H���� 3�#� g�����ʘ��(�h�G��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�#���"�p"  ����F�P3�3�d� �4Μ�)�r��)�r��)P| ͑�3Bp8^���eK�Ȋ���@&FrV_�1�0��e��C(�&bFa3����d^DU���eBp8^�М3S��9NS��9NS��*��$h&��8�B�� g�$*�S��$�_��`N$�2"PȉC"%��2"PȉC"%��2"PȉC"*����4#��pA9NS��A�eL���_����fY �k5�±|I$���A �2aD�	��������������������������������������������������������������������������������������������������������������������������������������$�2c�D�k5�J%�"���2d͉�6 x��)�r���7��xC �&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��@�Cs��C �R�`3� 2��q��Q�2NS��9NS��9NS�F�И��Nzd������q�Ȗ)�I�r��)�r��)�r��)�T 0X,f��h�g���e��Gdv��!�%�2d������������������������$�@B��)
�T*�LL@�L�2A(<�9NS��9NS��9NSdd��YU3M�D���6  2�O	�R'�<d���9NS��9NS��9NPygE8�>���� �pf�1�mrg�f��S���)�<�৒<B4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��<�G��#��د�>)�X3� 
��r�F p)�I�#L��r��)�r��)�r���ə��f K���\�ļ�����ac,eYxW�1 ��z+�,و�2NS��9NS��9NS��9M��3A���f��� 2�i>@T2V�Q,	Ē�DJ(dD���DJ(dD���DJ(dD���DX� �Z  �pA9NS��3L�4ʙS*
����2̲A��k5��d�H�$	�&$O�������������������������������������������������������������������������������������������������������������������������������������D�&L�2c�D�k5�J%�"���2d͉�6 l')�r��)�n2%����nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��*�@*q� �	�B|f� ,���#&f��)�r��)�r��(<�3�0Y���tF�Ӕ�9NS��9NS��9NP�|�i��`��3񟍀@�3�@�Pk5�������������������������񁁀P(lM��3񟍀	@�W*�d%�)�r��)�r��)�|�I	��<M��0�|�)�r��)�r��)�r���: ��20�fD^e\S"�
�\��S���)�<�৒<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��<�G��5S&�C2�� �3�*s$F���:r��)�r��)�r��)P| �М3f�@�͘��16b�34�> g)�r��)�r��)�r����p�7�g�Q�)V�	S�����P2�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��*���	P| �S��3L�4ʙS*
�����b��k5�I !���dɄ	$H@�?�����������������������������������������������������������������������������������������������������������������������������������@�< H��"I�&000Q(�Mf�YD�Q&L����&L��6&����9NR����)
J�@@T2���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ�� ���ĩr0�A6O��� 	�R�34�9NS��9NS��9NS��9NS��9NS��9L�4� �0�~?��3&dP(��H��������������������������2`�:��/G����?�P
 EAPg�)�r��)�r��)�r��)�r��)�r��(<�3�1~	J��Ɂ���3? �� 3�E
�D�eL!<�৒<B4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�S@��S�
!#���"�p"G� �L�����q�|��:r��)�r��)�r��)�r��)�r��)�r��)�r�#&f�ʨ��,_�8@e� � � �B0J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD��@�F )V�<NS��9EAPgS*eA@�W����Y�H5��b��_I #,�H&L�@�?�������������������������������������������������������������������������������������������������������������������������������������dɓ&L�IJ%Y��Q(�I�'���̲A ؛b �&�r��)�r��)
J�@@T2���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɰ��2�*�zM��'��)
��(<�9NS��9NS��9NS��9NS����`�ŋ @��8d�zAА000$O��������������������������L�2�D�(
��讙���X,�9NS��9NS��9NS��9NS��9NQN2O�)# 0H)��@�!�@C&�P!�0�h�G��F�D#@��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��D#@��Q�(�hB4
`h�eLxB�ey�p73�f8�N	��J#L��r��)�r��)�r��)�r��)�r��)� �pA3M�D&�r��x��PP����'X�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC",	ĀR�x8 ��)�r��i�eL���_����
±|k5��$��H$&L H���������������������������������������������������������������������������������������������������������������������������������������&L�2d��,�Q(��f�XV/��'���ɓ&lM�� @a9NS��9FqSa����@� ��y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���T�R/FzB� � *�&�ə�)�r��)�r��)�r��)�r�a!��3��6&�B@���2d������������������������������Y �k5�͉�6&TʙS4�3NS��9NS��9NS��9NS��9NS�F���Bq�� W� h^@�T�u�{<�৒<�G��H�S�
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x)�04
y#�L��S�W��L�O�����)�r��)�r��)�r��)�r��)P| ͑�0YU6e�� �'�i>@�@�U!,	Ē�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8�
U���9NQPT�TʙPP(���������k5��d�H```�2aD�	��������������������������������������������������������������������������������������������������������������������������������������&L�2d�
%���k�b��2����2f@��ŋ�)�r��8����h��"�ds����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��a"�1�L�BHU#4�dM��3NS��9NS��9NS��9NS���r2@� dЬ_�ɓ���������������������������$�Q(�F�؛�2�Q�� �@�����9NS��9NS��9NS��9NS��9E8�>�*�0��>GQL��
y#�O$x)���F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��D#@��<�G��H�R:�`����� h^ ϠpA #>r��)�r��)�r��)�r��)� �pA3M�D&�r��x�J�'	(W�|X�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2#9�W�*���	P| �S��A�eL���_�����f�Y��I$��	�&$O'������������������������������������������������������������������������������������������������������������������������������������ H��"I�&000Q(�Mf�X�+�ɓ����ɓ
�9NS��9Bq�� �Z  � ��y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s�������� N �'�eTD�9NS��9NS��9NS��9A`�X ��?���2���/F�Y��2��������������������������"L�A BA�2��8@� 6!�0�*��9NS��9NS��9NS��9NS��9NS�&/�(�!80�3(`E
�D���/b�S�
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
y#�D#@�u�{�'��\@��x�9~# 8�$�9NS��9NS��9NS��9M��0�e!M�b�&�	�*�z7<J�d#�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2#9�W�*���	�r��)�f��TʙPP(������b��k5�I "dɓ&L H���������������������������������������������������������������������������������������������������������������������������������������$�2c�D�k5���L�?���L�1@�PX�c��9NS�'HS=	!T�T2���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��#4�&i�ȟ �r��)�r��)�r��)�r��(<�3�\���H��g�`blA@�Q�H$������������������������2f�Y�P("�T�LLK,@(�A�r��)�r��)�r��)�r���9NS��9NS��9NPygBb��9� �3�/2�xB�j2�04
y#�O$x)��S@��L�F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S�
y#�O$x)��SP!�1�mrT0����� F|S����9NS��9NS��9NS��> `�pA3M�D������1*@�$�_��`N$�2"PȉC",	Ē�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dFr)���
U���9NS4�3L��2��P+����,�$�f�XV/�$����2d��'�������������������������������������������������������������������������������������������������������������������������������������	L�2dɌ
±|k5����V&L����&L�I���,X�9NS���Q�!> �����s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��:P2�%N "����3NS��9NS��9NS��9NS��9NR����0LX�b�/��#�;@P(001����������������������2d�%�a�sblM��C(�?�њf��h<�3�)�r��)�r��)�r���P_�|�#8X�3������T����)�r��)�r��(�'��X�ɳ2��ʹ��˓>�4��)�<���Q�(�h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!��F�O$x)�04
GQL�_|`E�	�� W���=2`�g>#L��r��)�r��)�r��)�|�HN2��p��*b��:P2Ȧb�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��E3�J�@A���r��)�*
�8ʙS*
�����b��k5�I !���dɄ	�������������������������������������������������������������������������������������������������������������������������������������&L�2d�
%���k/��X�H2����@�"�@��b�)�r��(N2��zB� "�ds����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<J�@E '�#86g)�r��)��!P���`�dr��)�r��)�r��(<�2D|��xbbb*�P��	$�@�?�������������������L�2I$�� ��G�2�Tʁ�xd�����g)�r��)�r��)�r��A�	O�pɑ��3�/�>e e�4S1p�����d� J�A~*��r��)�r��)�#L�<�3��H)��x`E���>GQL�@��<B4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
!��H�S@�u�{rg�f�&�C2�� �3	�\���4Μ�)�r��)�r��)�r��)��π�e!@)V�(q%�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��E3�J�@A���T 3��9L�4�2�Tʂ�@����̳,�k5��b��$�@FY �L�2d��������������������������������������������������������������������������������������������������������������������������������������$H@�$ɓ�b�BA|_
ĂA������(
 �$	����9NS�UDD`��*�@�e!���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8�� O6Fpl�S��9NQN0�0S��2��6eTT��4�9NS��9NS��9BPy�d�����<�H� ��H H�������������������	L�2�D�P(ə3 `���F�!�1�f���4Μ�)�r��)�r��)�T 3�/�0��6��$|�h0'
F����"�n �hUJ�3A�8�l��� ���1	O�p�> g)�r��)�r��)�#L� F|�h� }�x@�W��#��؄h��)���04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!��F�H�)��+�O�,��3� 
��r�F p)�I�#L��r��)�r��)�r��)�r��)�l��ٕq���e!`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��*���	�r��(�*�*eL�(
����```V��Y��I$��	�&$O'������������������������������������������������������������������������������������������������������������������������������������ H�dɓ&L```�/�cY��_± �e����P( H��t�9NR���ʨ��l� EP��ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8�� O6Fpl�S��9NP8�":h�9��K�e����T�����͐<�3�)�r��)�r��)�f��h��TʙR8G�@�P$��AD����������������ɓ&I �C��T*������~? `d�����t�9NS��9NS��9NR�����>
�����M���P8
 J�T�=9���F�z4sѣ���hUJ�3A�9x�����2�)��)�r��)�r��)�#L�L_�R�=2``�`��fz�\��S���)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��C*c��(�̫��F���� ��<�3�)�r��)�r��)�r��)�r��)�r����"^ Џ�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'J�@A���T 3��9L�4�2�Tʂ�@����̳,�k5��b��(�J&Y �L�0�"B��������������������������������������������������������������������������������������������������������������������������������������D�&L�2c�D�k5��f�d������"J���~	A���r��(,���&�	�a"�&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��F%H�� l��ٜ�)�r�����G�g�:@Yb���*�>��@hȕp�D� ���t�9NS��9NS��9EAPg `?���#��@�V/���"���������������"I$��``lM��>�O�TʙP6�&	�`�Y�r��)�r��)�r��)P| ��ૄ�x�����R F^T�d��	U*��G=9���F�z4sѣ���h�G=9���F��"�T�d���f
�S� S����eA�9NS��9NS��9NS�&/�(�!80�2��ʹ���ʘB4
!��F�D#@��Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��Q�(�hB4
`h��)�<�৒<���/`���=>������ �,L�g�S��9NS��9NS��9J��l��ٙ�U	(���6b�> g)�r��(N2��`3�`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȊ�d# �D')�r����3���2��P+���񁁃Y��k5��$��H$&L H���������������������������������������������������������������������������������������������������������������������������������������$�2c�D�k5��f�A �����D�
����σ��9NPx8 ��(�A���ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��@�B�@	�����r��(l�2���*�X���� ,�e� U��Ч��HT#�0ygNS��9NS��9NS��a!����#�p$�LMf�Y2d�������������@�# �:�A�3&d��ıb�\���X,r��)�r��)�r��)�T 0���^�8,��9�	 �3A�9��R��z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�AРpe e�p��~2g�J�A~9NS��9NS��9NS�S���� �,�9~2��ʹ����>`hB4
!��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!04
!<���R:�`���3�3E2+ ��@���F����d��ygNS��9NS��9NS��9M��3Af�@�"��	���2�Q���	��W71�1r��)�T 0�e!H�g���I(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���@)V�<NS��9L�4�2�Tʂ�@�����f�Y��k$�@FY �L�2d��������������������������������������������������������������������������������������������������������������������������������������$I2dɓ&000_°:��Y��H$�����?���X,�9NS�UDD`��*�@7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���P Bx��3�fr��)��π�0 
��� ,�e�,@Yb�X\r:h� ���	��&2`0Y�9NS��9NS��9NPX,Uʹ� He��d�z5��cD������������&L�|_
��!�P�F~3�����b��3�Py�r��)�r��)�r��)P| ς����Fp��"	�3#,��J���M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�S`�d p���  �g�P_���r��)�r��)�r���d��H)��xS"�
+�O��S���(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!��5S(W$x@�@� �pe$d� ygNS��9NS��9NS��>�$l���/fT��������ВO���A� ����¼ ��)�r��'HQh!�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'J�@A���T 3��9L�4�2�Tʂ�@����$H�����k5��d�H```�2aD��"������������������������������������������������������������������������������������������������������������������������������������2dɓ&000Q(�Mf�Y��k$��"����)
G�����)�r���A6O�"�ds����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<Hĩp���3��9NP,�����H,@Yb�X���� ,�e�, �WH�U�x2����f
p�Ʉ����9NS��9NS��9A`�XLÎ9�blA�t$&L H��������� H��"F@�Q�6&��}>����3@��2@�X,�9NS��9NS��9NS��> a)��x6c$ ��� �z*r2^P��L�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"� �R���`Ng�HWј*����P_�S��9NS��9NS���$�*�H�20� }�	�证>GQL��(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��S�
y#�D#@�u�{5S мD^e\��ٕ9�	��J#L��r��)�r��)�r��)� �f L�xb�U�g/`#��C3�3 ���H�����q��\ ��PgT$���9NS�UDH�g���I(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD��@�F )V�<NS��9EAPgS*eA@�W����ɓ5��b��_I #,�H&L�@�!D��������������������������������������������������������������������������������������������������������������������������������������"I�&L�1����D��� �k5�	_���␤)���X,r��)�8@e�7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<@�@�nx<�8�� O6Fpl�S��9BPy��W���� ,�e�,@Yb�X���� ,�����U�x2��,lʨ��#��9NS��9NS����a0L8�&&"�U
�P(001�������$�$�t$ ^��#�q�0� �3�S��9NS��9NS��9J��|�ɑ��3�3Epe e�4�%T�f���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9����L���yD	 aNl�,� �P| �S��9NS��9NS�F�И�����0�0̠!��"GQL�@��Q�(�hB4
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�(�h�G��H�S@�u�{P�D3� 3��������'�<�3�)�r��)�r��)�T 2����8f��_�x�@ D'��3��WBHy3�3	��\~>������q��\~>� &��_�S��9NPYU6�`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȌ�S1_��D!(<�9NS��3L�*eL�(
�����2��Y��k5�I #,�H&L�@�?��������������������������������������������������������������������������������������������������������������������������������������"I�&000_°:��Y��H$aD�������?��`���9NPx8 �q��6�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��S�� ��dg��9NS�6@``@q�,@Yb�X���� ,�e�,@Yb�@g��e��
�y%�	V ��=�1�F��)�r��)�r��)�d��� @a111*EH��$�@_�����&L���k
H�"�/��?����i�r��)�r��)�r��)�r�A~�����0�6 �l����!
F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�NFK�^`�A�9�8,�|�%A�9NS��9NS��9NPygBb��9�s96fQ�W<�x5S<���Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x)�<��u�{�'��\@�D^e\�9~D's$F���:r��)�r��)�r��)�l���6bf���V�/3�s��2��f!�f����}.?K��������}.?K����p0	��z+�P| �S��*�N2��`3�`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȌ�S1_��D')�r����3���2��P+���񁁁XV/�f�Y$�&L�@�!D�	������������������������������������������������������������������������������������������������������������������������������������	��&L�2d���V5��`�:?�������,9NS����	Wpla�f�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8�� O6Fpl�S��9@`�d�3�@�e�,@Yb�X���� ,�e�,@Yb�X����/32U䗐l%��2�,	�>g�8d�h<F�Ӕ�9NS��9NS��3L�4���2fJ�D�Q&L����&L�D�Q1Gdv�����?�њf��hJ>S��9NS��9NS��9O�����Bp<��P �~	�p�9/(UJ�9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSB��Q��������ɟ�a(|��> g)�r��)�r��)�)�I�F p�D^e\S"�
+�O���F�D#@��L�04
`h��)��S@��L�04
`h��)�<�৒<��)�ʘ�6���0��AL��H�S����9NS��9NS��9NS����Y�%��W�nb"�DF&G3 �J��f!�f����}.?K��������}.?K��������}.?K���&�xc�2NS��9Bq��# A�q$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���Dg"��� �Z  �pA9NS���8�*eL�(
�����2��Y�V��I$e�	ɓ'��������������������������������������������������������������������������������������������������������������������������������������"B�&L����D�Q5��`�:?�������,9NS��> `�pA*�.�l#<��y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��1*@� ��dg��9NS�F���1��H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd��g�:X�,2��#�z3�H&���i�9NS��9NS��9BPy���02�Tʙ�2fJ�D�Q&L���&L�I��H
p��  	��">d�`�XJ>S��9NS��9NS��*�J|�L�/e�ɟʹ�m/0W#4�%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"� �R���L2ٙ�f2@ ��1>
��T 3��9NS��9NS�F��ygD3��S83� 
�"���_|���/b�Q�(�h��)��S@��L�04
`h��)�<�৒<��)E0^�|	�!L��)�� W���M�S��0����4Μ�)�r��)�r��)�T 24'�Y�&H���g"��	�ٜ����C(�&bFa?K��������}.?K��������}.?K��������}.?K���&�xb����)�T 0YU# A�q$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���Dg"��� �Z  �pA*��r��i�f�S*eA@�W������_�f�I$e�	ɓ'��������������������������������������������������������������������������������������������������������������������������������������"I�&L�1�������t$�f�����"���:��*eL�,9NS����	Wpl1*@���y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<@�@�T�( !<@���9NS��	A��Xφy�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@ 
����L� ��&h�G�a(<�9NS��9NS��9NS4�3@('����}>��X�/��&000+��P(*EH����8�Cc4�3BPy�r��)�r��)�r��)P| ς�� �PS���S� @��	#4���qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qS@�U1�	���
�3@0��t%> ���)�r��)�r���4΃��:����B���� 3�E
�D���/b�S�
!��F�L���H�Q�(�h��)�ʘ͢ �ef@�3�d� �4Μ�)�r��)�r��)�T 1�a�+�	W71c(����&䬿�bFa3�3	��\~>������q��\~>������q��\~>������q��\~>�����`H���')�r��8�B��A�'J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8�
U���9NQPT�TʙPP(���������k5��d�H```�2aD���������������������������������������������������������������������������������������������������������������������������������������&L����D�Q5��f�Y�``c����t	A�r��)�2�g#�	���s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q � l��ٜ�)�r��f�,g�<���X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]W��Z�?�$df�h�	��<�3�)�r��)�r��)���('���e��*�P�*EH�����?����">d�`�Y�r��)�r��)�r��)P| ��૊����M���S���%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѠ	U*�����I���P� �P| �S��9NS��9NS�F�Үd���Bpa�fP����E0^�#@��<B4
!��H�Q�)E0^�|	� E�&~^?�_���Ʉ��%��t�9NS��9NS��9NS��34'��f���Ȋ�{ ���Y��2��	� �?K��������}.?K��������}.?K��������}.?K��������}.?K����p0	�$^ ������9BPy�*�%��`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȌ�S1_��D%A�9NS�Tq�2�T
���000k5��f�Y$�&L�@�!D�	������������������������������������������������������������������������������������������������������������������������������������$I2dɓ&000Q(�Mf�Y��k����BAAPg�)�r����=2�F%H��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��F%H�� l��ٜ�)�r�����G�g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,�f*�:h*ȫb�G8Ld�Py�r��)�r��)�r��0Y��C�x��xL��X,�9NS��9NS��9NS��> a)��x6c$ ���R F^T�d��	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aҧ#%�2�2�f�K�?���J��r��)�r��)�r��(L_�R�=2`ng&��"�*�ɴD�eL!<���M@�Tǀ4/�@���F�F����8�>S��9NS��9NS��9J��6b���UJ��,eXg�A�����C(�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q���/ l|�I�r��(,����4#Ł8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"3�L�~�R�x8 ��)�r��i�eL���_��� H����Y��+
��$�2̲A2d��������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000_°:��t	�H����t	A�r��)�F�h8��9� Nnx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d*q � l��ٜ�)�r��f�,g�<���X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��U�t*�<U�V�	��6eTT��4�9NS��9NS��9J��r��)�r��)�r��)�r���8d���)�`l)̀g�HWњ	�Q��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4(Hx/�>_���ɑ���*��r��)�r��)�r���d�`g���E�U�2+ �ɴD`E�	�� W���=2`�g>r��)�r��)�r��)�T 1�`��p��R�2"�^�&Gc��f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����p0	�$^ ب> g)�r����"J�@Kq$���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���Dg"��� �Z  �pA9NS��3L�4ʙS*
����&L���k5��d�H�$	�&$H@�?������������������������������������������������������������������������������������������������������������������������������������ H�dɓ&L```�/�cY���� �I����� �i�f��)�r����=2�F%H��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��T�( !<@���9NS��	A��X\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�|3�*�#�fz88lʨ��#��9NS��9NS��9NS��9NS��9O�����E@yT�P&�̌�L2�pn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���%T�c,�A6fdٌ� d���|��> g)�r��)�r��)�#L� F|��B��r�d`!P��"4F��ygNS��9NS��9NS��6FL��1_�E# 	�X�0�s1�rV_�����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K���&�xc�2NS��9AeTD�h��Ȧb�IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��E3�J�@A���r��)�*
�8ʙS*
����2̲@�+ƳY��Id�A2d��������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000_±��k5��d�H����Y�� ���4�9NS��#A4	�ze�J�'7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���P Bx��3�fr��)�� �0 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb����φy���2�`cfUE@,���:r��)�r��)�r��)�r��(J|��ɟ��~	�p�����L�A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�a*������L���g��x	O�p�> g)�r��)�r��)�#L�'�<�3�)�r��)�r��)�r���34'��f���Ȋ���@&FrV_�1�0�ϸ���\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q���$^ ب> g)�r���pA �Z &r)���PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"3�L�~�R�x8 ���9NS4�3L��2��P+����	L�1XV/�b��$�@Cɓ&L�������������������������������������������������������������������������������������������������������������������������������������@�< H��"I�&000Q(�A�t$��H$�@_�����f�4�3NS��9M��0�g�Q�ĩss����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y�e!� N Bx��3�fr��)�� �1��H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���P�$@Yb� "�>��3���W#�z3�H&��S��9NS��9NS��9NS��`p�������z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�%T�eNFK� H�!
s`�`��S��9NS��9NS��9NS��9NS��9NR���͘�/Ǣ��R�9{ ����P3���������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��Y�a������9NPYU �Z &r)���PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"*��� R�x8 ��)�r����2�Tʂ�@����̳,�+
���k$�@Cɓ'�	��������������������������������������������������������������������������������������������������������������������������������������&L����|_
ƳY�BA$�'������|bbbd���9NS��6FL� !<@���f�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8�� O6Fpl�S��9A�i� ��� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����29�&rg�<��HR�*b:R23A4T#�0ygNS��9NS��9NS��	O�pg ���� �z
C���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4���yK���� �ϛ!�9NS��9NS��9NS��9NS��*�ϊ�0��/fT������|��Y��2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>���Ø�3����<d��)�r�ʨ�*�,	Ē�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�h�����> g)�r��i�eL���_����&LV��X�/�%��H$&L H��"�������������������������������������������������������������������������������������������������������������������������������������$�2dɓ(�J&�Y�BA$�'������|bbbd���9NS��6FL� !<@��Pnx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d#�	�O6Fpl�S��9@`�dg���|3� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yc#��g �*�@hS��FFh&��qr��)�r��)�r��)P| ��૊pX�4WR F^T�d�����z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �hP8
�0�6 % �S��9NS��9NS��9NS��6FL��1d��R�8�/����(�e��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.�1�F�>�$�9NR������h���IC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��B0J�@A���r��)�*
�8ʙS*
����&L���k5��d�H�$	�&$O��������������������������������������������������������������������������������������������������������������������������������������2dɓ(�J&�Y�BA$�����k5����">d�S��9M��3@O*q�&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��T�( !<@���9NS���͐Xφy�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb��9W��X���M��t�9NS��9NS��9NS��> a)��`aNl�3rT�d�����z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A���Lf�s) #/��'��?��P�> g)�r��)�r��)�r���<d����^ Ex�@ D'���@ #9+/���Q�O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.�1�F�>�$�9NS�UD@)V�	`N$�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq �D �4Μ�)�f��i�2�T
���L�3Y��k5��$��H$&L�2������������������������������������������������������������������������������������������������������������������������������������D�L�2dɌ���� BA$�'����J%�/��2D|��)�r�#&f��� *q�&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��T�( !<@���9NS��	A��X\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y`@qʘ��TT#�3��9NS��9NS��9NS��*�J|�8@�1$|�����*�S7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M6�_�)���!_F`�p<���8T 3��9NS��9NS��9NS��34g
�UJ���dv9�fbFa3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\9�`�{2��<d��)�r�ʨ�����E�8�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"3�L�~�R�x8 ��)�r��i�eL���_��� H�dɚ�f�Y��I$��	�&$O'������������������������������������������������������������������������������������������������������������������������������������D�	$I2d���V5��`�:	$�@�?��������	�`��9NS�����~ ��`�7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s��J�' !<@���9NS���͐X\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�L�x�1�9NS��9NS��9NS��9NS��*�J|�L�/c0T �ٙ��	��U1�F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qS@�U2�#%�/0W ���0�>
��T 3��9NS��9NS��9NS��*�~=�e��ВL�2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\9�c0��|�I�r��(<���	����EP2�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"3�L�~�R�x8 ��)�r����2�Tʂ�@�����
%���k$�@FY �L�0�"B��������������������������������������������������������������������������������������������������������������������������������������D�&L�2c�|+�f�t	� H����I �P�A0L�)�r� �3� ��Pnx<��2����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s�����bT�8	�����r��(l��ppφy�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���G3�@�/�&2g)�r��)�r��)�r��)�r��)�r�A~	��:l�H M����	U/��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��A�� �323@�PF�\�> g)�r��)�r��)�r��)�r��(,و�2"�g%e�?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K�����Cٕ>�$�9NS���pA6O�@�F	C"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��E3�J�@A���r��)�f��i�2�T
���L�1XV/�f�Y$�2��dɄ	�������������������������������������������������������������������������������������������������������������������������������������&L�2d�
%���kAАI ������e���1�r��)�#0� 
�@E�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8�� O6Fpl�S��9@`�d�3�@�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,����3��28)�c&r��)�r���: ��*s�&e$d��F�Ӕ�9NS��9NS��>
��	@3f2@ �l����!
F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��a*������L�����ɟ�a(|��9NS��9NS��9NS��9NS��9NR�����_���>L�2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>���Ø��*|�I�r��(<D`��T�`�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȌ�S1_��D%A�9NS��3L�*eL�(
�����2b��_�f�I$000L�0�"B�'������������������������������������������������������������������������������������������������������������������������������������ H��"I�&000_±��k�E�D H����I �P�A0L�)�r� �3� ��Pnx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��S�� ��dg��9NS�F���0 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt�R�)�c&r��)�r� g���M��E�U������i��<�3�)�r��)�r��)P| ʃ�	@2�d��p���8^���Q��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4�AРp"�ٙ��* @N�Д�
��r��)�r��)�r��)�r��)�r��)�r����66��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K�����Cٕ6FL�9NS��#A43ВH�B0J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dFr)���
U���9NQPT�TʙPP(�����2̲@�+°�_I #,�H&L�@�?�������������������������������������������������������������������������������������������������������������������������������������	L�2dɌ��k5���t$@@ �"���$�C(er�FNS��9O�x��� ^��	3s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y�e!S�� ��dg��9NS�F���0 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt�R�)�c&r��)�r�"�\�U>M�'ɴD`E�	�� W���M�S��0����4Μ�)�r��)�r��A�*�ϛ!S�����2�2�pn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѠ	U*�����0�6 ���ϛ!�*�P| �S��9NS��9NS�F��PT�0L `�`L��4Μ�)�r��)P| ̑xca �L��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3������ʟA~9NS��#A43ВH�B0J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dFr)�����x!(<�9NS��3L�*eL�(
�����2b��_�f�I$e�	ɓ'������������������������������������������������������������������������������������������������������������������������������������ H�$H@�$ɓ/��X�k5���H(�J!D���񁁃���!�0�9NS��*��,_�*�z EP��ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��(
�@E '�#86g)�r��0Y�3���>��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ҭ28)�c&r��)�r�TL�A�"��G6�� м,��2��ʸa�8�N	��J#L��r��)�r��)�r��g͐�3�e��9����S���"�9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSJ�����@���~	�f2@�#K�J|�A�9NS��9NS��9NS�%�i�f��xeL��>�O��U
�T*�P�C(q�A�r��)�r����66��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K�����Cٕ6FL�9NS����	����EP2�PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC",	ė�4#���"r��)�*
�8ʙS*
����&L���k5��d�H```�2aD�������������������������������������������������������������������������������������������������������������������������������������$I2dɓ&000Q(�Mf�X(
/��X H����000}>�D0��)�r���<d���"T�R/F�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��R�'�#86g)�r��(<� � ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �W@�/�&2g)�r���4ΙT3(c��"��G6��(W �����"���(�̫��F�P3�3��4Μ�)�r��)�r��)P| ��ૌ�`aNlG����yM�M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�%T�c4S3=2B��
s`
pX �P�*��r��)�r��)�r��(, �@�����/��*EH�
�D�e�	 �:ə3 l �X,�9NS��> fH����@&G��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��Y���eM��3NS��9H�M�$�R*����DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�x�Q����)�*
�8ʙS*
����&L���k5��d�H```�2aD�	$O������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�/�cY���� �/�`�"������#�pCar��)��σ4�dFi>M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q � l��ٜ�)�r��f�,�9e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,����3�:eK��	���r��)�d`!P̠!��h�#�DA�"����"|�DO�h��mȬ���fAL�A #>)�I�r��)�r��)�r��(J|�8+�g�>$f�p��Lsѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aҧ#%�2�2�8_�|ٌ� ��t%> ���)�r��)�r��)���`�& @a2�TʟO�� d�:��,�H'��f�X�C(&	�c��9NR���"��� ������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\g%e�ٕ6FL�9NS�����l�*����DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�x�Q����)�f��i�2�T
����"I�&k5��f�Y$�2̲A2d����������������������������������������������������������������������������������������������������������������������������������������&L�2c�DB@(
/��X H����000G��C�)�r� �f���SH��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d7<J�@E '�#86g)�r��(<� � ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,ds0L���p�ɜ�)�r���:d`!P̠!��h�#�DA�"����"|�DO�h��msh��mȬ��0��AL�A #>)�I�r��)�r��)�r��)�T�&F���*�=2B���aL��U1�F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ������	�	 �)̀3�e�|�%A�9NS��9NS��9NS�%� �X,�Q	@��
�T*�!HR$�@AD���```��� 09NS��*��/ ll 	���\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>���Ø��*F��r��)��!>X�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��I�*�')�r��i�f�S*eA@�W�����D�k5�I #,�H&L�@�!D��������������������������������������������������������������������������������������������������������������������������������������"I�&L�2A �(�J&�Y�
��$O���#�p� P
 NS��9BPy�f����#�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%N "����3��9NP,�����H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@2��S��L�9NS��20�fP�ɴD͢'ɴD�6��&���"|�DO�h�#�DA�"|�DO�h�����fz }���񔑐�'�<�3�)�r��)�r��)P| ς�� �Pٌ�  �323A�3 J�T��M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�n �iS���Hx/�>l�H 2di{	O�p�> g)�r��)�r��)�r��`��&	��<2�Tʑ�8G�A��k&L����&L��6&����9NS�������~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q����/fT�34�9NS�)����U!%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��I�*�%A�9NS�Tq�2�T
���L�1XV/�f�Y$�2��dɄ	�������������������������������������������������������������������������������������������������������������������������������������@�$ɓ&L����D�Q5��`�P(�/�`�"������#�p �3��9NS��70���y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<@�@�T�( !<@���9NS���͐X\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�3%PL�x�1�9NS����t��B�!�@C&�G6��&���"|�DO�h��m>M�'ɴD�6��&�G6��(W'ɴDS"�
  ����x�9~# 8�$���t�9NS��9NS��9O��� �Pٌ� �O�����J���M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�@�(e�a���� ���,3��A>
��T 3��9NS��9NS��	A���*�
D	��~C(e�� a�rHL�?����&L��2����9NS����^�&G`��p	����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3������ʛ#&f��)�r�#86`p��20��C"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'^ Џʨ��r��)�f��TʙPP(�����2̲@�+±|_I !���dɓ&O��������������������������������������������������������������������������������������������������������������������������������������"B�&L����D�Q5��`�P(�/�`�"���2d�ə3 ���:r��)P| ��q�# A���s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y#�	�O6Fpl�S��9BPy��W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���T�*^8Ld�S��9A�i�20�fP�ɴD͢ �m>M�'ɴD�6��&���"|�DO�h��m>M� �msh�"�p"����< zg�@�73�fT�L&/�(<�3�)�r��)�r��)�T 1�6B���/�>e e�@�(�A��F�z4sѣ���h�G=9���F�z4sѣ���hUJ�T�d��R F^U��i~2g�&F����
��r��)�r��)�r��(<�3�0L  	���0g�2fLȠP(5��fY ��������"L��/@x��)�r�����^�&Gg��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��Y�a��34�9NS�����QT�`�2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq$`3�,�����9NQPT�TʙPP(����2d�f�Y��k$�@Cɓ'�	������������������������������������������������������������������������������������������������������������������������������������	��$�2c��_��H�F�Y� H����000fLə �0�9NS��3M�D�x7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���P Bx��3�fr��)��#=3�@�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����T�
p�ɜ�)�r�����C2��<�xsh�#�DA�"|�DO�h��m>M�'ɴD�6��&���"��G6��9�D͢ ���"�p"|�DH���p F@��M��!8��"4F�Ӕ�9NS��9NS��*�ϛ!S���S� �@�ʜ����A��F�z4sѣ���h�G=9��qSB��P��A6fd ���,F�\�> g)�r��)�r��)�r��H��  �����lT*�P�)
D�H H�������$H�P( @a��t�9NR����U	(/3��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/����8f�)�r�#86`p��*����DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�x�Q��9NS4�3L��2��P+����dɊ±|+��D�Q2��dɄ	$O������������������������������������������������������������������������������������������������������������������������������������$�2dɓ$�@E�D�k5��@�Y��L�?���L�2�T����)�r��)�n2$`3����nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%N "����3��9NP,� e�� U� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����/32U tʗ�N3��9NPygL�*�1�msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh��mXqey�p0�0q���F�Ӕ�9NS��9NS��*�J|�8XS� ��\�9/(UJ�n �h�G=n �hUJ�3A�9����s4�_����g�P_�S��9NS��9NS��9EAPga!��H fLə
�|+&O���������
�8<�3�)�r�����^�&Gg��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��Yʹ���2fi�r��)�3�f�#��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq$`3�,����)�r����2�Tʂ�@����ɓ&k5��f�Y$�2��dɄ	�������������������������������������������������������������������������������������������������������������������������������������$�2c�DB@(
5��dɓ����ɓ6&�ؖ,X�> g)�r��8����� EP� t�d7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<J�@E '�#86g)�r��0Y� � ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� �/�&2g)�r���4ΙT3(c��"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"����"|�DO h^\@��0a�U4T@σ��:#L��r��)�r��)�T 0��p<��b H���)�S���9/(��!M����	��:� �P| �S��9NS��9NS����fi�f�`~?�P�F�؛P(000L�?�������� H�@�P8ㄠ���9NS����^�&Gg��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��Yʹ���2fi�r��)�3�f�#��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq$`3�,����)�r��i�eL���_����&L�k5��f�I$e�	ɓ&L��������������������������������������������������������������������������������������������������������������������������������������D�	L�1����D��� 
�f��"���@�"��`�Y�r��(,����(�J�'�e!���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��(ĩp���3��9NPyg@2��|3� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�tʗ�N3��9NS���B�!�@C&�G6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h�#�DA+���"�"�̠!� Ϡp
g�ygNS��9NS��9NS��> g�P_��^�8,��� �d��,	@3�/�A�9NS��9NS��9NP�|�`��&	��LLLJ�R*B�@��k5�d�G���������$P(  	������9NS��
�IE�dv	� �?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/�W71#Bp�9NS��6Fpl�`�����J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8�0�UDBPy�r��(�*�*eL�(
����D�&L�k5��f�I$000L�0�"x@�?������������������������������������������������������������������������������������������������������������������������������������D�	L�1������f�X(
5��aD����I$���#����9NSdg��7��x�J�'7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<J�@E '�#86g)�r���4΀e���g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� �/�&2g)�r���4ΙT3(c��"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh�#�DA+�E
�D�6��dVA����+���񔑐�'��r��)�r��)�r��A�>
��T 2����)�r��)�r��)�#L�f��x�������lM���
%������������	(
 �J��r��)P| �p� %�dv	� �?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/�W71#Bp�9NS��6Fpl���d`5�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$�x�Q����)�*
�8ʙS*
����(�J&�Y��Id�A2d��'�������������������������������������������������������������������������������������������������������������������������������������	$I2d�
%�:��P(k5�ɓ'����@�%�@�H��#��9NR4A�fX��zB�1T�Ѱ�y@�@�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��2����P Bx��3�fr��)��#=3�@�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����T�
p�ɜ�)�r��F��6��9�D͢'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� ����mȬ�&g�~^?�_���b���)�r��)�r��)�r��)�r��)�r��(,�C,X���̙�2(

%�2d�������������"E�@��σ��9NQ�+�	{ ���e��}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K�䬿�\�č	�0�9NS�����Q���J(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ(dE�8���xUDNS��9L�4�2�Tʂ�@����ɓ&+
���k$�@FY �L�0�"��������������������������������������������������������������������������������������������������������������������������������������D�&L�2d�H�Q(��f�P(k5�ɓ'����6&�؟���$G̑�r��)�2fhN2��0�L��R��f0I�!�C �2����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���@	�����r��(J> 2���*�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yc`� #��*�:eK��	���r��)�d`!P̠!� h^�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DA�"����"|�DO h^��韁 W���0������4Μ�)�r��)�r��)�r��)�r��`�$G̐������}>�blA�t$d�@@�?������������D��ŋ����9NR����^ K����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/�U*�3��8f�)�r�#&f�q��20��C"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%���(��I
���9NS$G̑�����k�����2���_
±|I$��	�&$H@�!D�������������������������������������������������������������������������������������������������������������������������������������	$I2d�
%���kAАk5�ɓ'������D�"� �&�#L��r��(J>��0�e!@O3ВH���^��g���&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��F%H�� l��ٜ�)�r��f�,�9e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����T�
p�ɜ�)�r���:8�N3(c��"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6�� м,��2��ʸ�ɳ*s�&	�p3��4Μ�)�r��)�r��)�r����*�\���ºbbb@�3����D�2aD���������������$	@�X,�9NS�g
�^�&GfbFa?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/�W71#Bp�9NS��6FL�*�.�P����2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȍ���g�Qπx�9NS�� �0̙�2I$�����@�&Y�H�b��k5�I #,�H&L�@�?�������������������������������������������������������������������������������������������������������������������������������������dɓ&L�IJ%t	 �P(�k5�&O����e�	�!ϧ����X,�9NS��9J��l��ل�)
3� �BHU"�f0I�� EP��ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��2����P Bx��3�fr��)��π�0 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����fJ��R�)�c&r��)�r�T3(c��"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD͢ �msh��mXqey�p0�0��L��'��r��)�r��)�*
�8f��#*eL�#�p��
����������������$Ha�pH��i�9NS�%�8/e�dv~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q������`�М3S��9O�x�*�.�P����2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"���3���
��r��(�*�*eL�a�p�"���&L��+ƳY��Id�A2d��������������������������������������������������������������������������������������������������������������������������������������� H�dɓ&L�H2�%���k�# t	ɓ�����2b�@������4�3NS��9NS��9NR���#86a8�B��� M��LU"� �����:P2�&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%N "����3��9NP,�����H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�2��S��L�9NS�F���Bp!�@C м9�D͢'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �msh��mȬ��x
g1~	NS��9NS��2D|����T��@�P(�J$ɓ����������������!� H	A���r��A�¼ ��	����\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����rV_�U�g�P&9NS��6Fplʸ˃`�+�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"*����8|�2��6FL�9NS���º@�3�I$����@�$ɓ5��f�Y��I&L H��"������������������������������������������������������������������������������������������������������������������������������������@�$ɓ&L����|_
ƳY�B��t$&O����D�2�P��C�)�r��)�r��)�r��A�6Fpl�q����  �'�i>Hĩss����y7<M��s����y7<M��s����y7<M��s����y7<M��:P28�� O6Fpl�S��9@`�d�3�@�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����T�
p�ɜ�)�r��F��6��9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"�\�(W'�4/Q�WD'��:r��)�r��`����d�z$�@_�����������������"CC�@�$�σ��9NP���2�,�C(�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\g%e�*�Xq�c��9NS�2J�˃`�+�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��'d`5�R��Dٖ/�<S��)�*
�8�b�d̙��D������ɓ(�J&�Y��&L H�$O������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�H2���VAА!F �:	�'�����1?��`�dr��)�r��)�r��)�r��)�l�����(	�	�B|���^�ĩss������ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��S��&�sdg��9NS�%� ``@q�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�2��S��L�9NS��20�fP�ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh��E`0�	��Jr��)�r�P
 H�#��������������������(
 �$	����9NR���͘�c(���2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����rV_��EZ�P&9NS��6FL�*�.�P����2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%P2�:P28���$�R�� *�'�<d��)�r�r�FLLLJ�2d�����```�Q(��f�HL�2dɄ	�������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�/�cY��!F �:	�/����&LP(����9NS��9J��T 3��9NS��9NS��6FL��QfX��	�B|f���J�'7<@�@�nx<��&�ɹ��nx<��&�ɹ��nx<��&��S�� ��dg��9NS�6@``@q�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�2��S��L�9NS�F��#
��e|�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴDB�>M�&~^2�29NS����tq�6&�ؓ&O������������������1	@�,9NS��> `�f FX�0�1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��Q�D9hl�	�r��)�$d��@�BPȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��I���l �^R0ૌ�6�n2 �pA>�$%�)�r��)�#�H�?��8GC����ɓ&k5��f�Y$&L�@�!D��������������������������������������������������������������������������������������������������������������������������������������"I�&L�1������f�X�!��H&L����&L��P(� H�9NS��9HМ3p� !8/`�NT 3��9NS��9NS��> f�ə���"l��A6O�1T��� Nnx<��&�ɹ��nx<��&�ɹ��nx<��&��S�� ��dg��9NS�6Fz88g�<���X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�*ȫbS��L�9NS�F��#
��e|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&�E
�D�6��D^e\�H��9NS�F��H���/AD�����������������1?��`�Y�r��(,و�2�,�C(�'��q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\g%e�L�U�Y�')�r���ə�d��P����2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"��I`N$$�_��{3$�`���?  �e!H�M�x�9NS��9NS��	A���f��� @P(&O����	e�d��D�k5��$����2d����������������������������������������������������������������������������������������������������������������������������������������	L�1������f�X�!��H&L����$P(����9NS��34��6	�"	�"*�Xr�z+�,و����)�r��)�r��)�2fh,���2���Q�F%H�� t�d7<M��s����y7<M��:P28��a��G#A49NS���͐Xφy�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt)�A��9NS��20�fP�ɴD͢'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DA+���(�̫�I��)�r���# d�@�?�����������������!HR?���X,�9NR���͘�c(���2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����rV_��EZ�1r��)�|�Ip3��+�%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%P2�a"�4#�\e���q��Qdd�Ӕ�9NS��9NS��9NS���C��2�f�_����ɓ�b�V/��I$e�	ɓ&L��������������������������������������������������������������������������������������������������������������������������������������D�&L�2c�DB@�!��H����D�
����σ��9NPY�"	��� ��P9�f� ���ae\����6�1|�I�r��)�r��)�r�#&f�ʨ��,_��!>F �<�R�� ��y7<M��s����y7<Hĩp�g�Q��MS��9A�i� � ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,�f*���T#�3��9NPygL�*�1�msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m>M� �msh��m3� 
񔑐�r��(J>���2� H���������������������2�T��)�r��p����a`�3� ~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����rV_��EZ�1r��)�|�HL3�(�t�d%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"PȉC",	Ė�@�@�^��	3=	!T�O	�R�����t�9NS��9NS��9NS��9NS�Tq���!K����,�$�f�Y��I$��	�&$O'������������������������������������������������������������������������������������������������������������������������������������ H�dɓ&L```�Q(��f�HR�@�Q2d����@�%�@�?���:r��)�6b������Lb�!���L &�	��U*�3���_�f�@� �r��)�r��)�r���<d�ʨ��,_�8@e� �bT�8*�@�e!���nx<��$bT�9p3����)�r���:�W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��U�O��G�g)�r��)���@C2��>M� �m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD͢ �msh�"�p"xB�ey�s)# 3��9NR������ d�@�?�����������������!HR?��⠨3�S��9Af�@���afbFa?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/��g"����)�r��f�&�p:P2�DJ(dD���DJ(dD���DJ(dD���DJ(dD���DJ`N$��j6B/)��4�dA���|�I�r��)�r��)�r��)�r��)�r���X,�?������D�&L�Q(���|Q(�L�A �2aD�	������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L```�Q(��f�B0�D�A������1?��Py�r��)�6b����&b�!�b�!�bg�@�/��
�V���6�1|�I�r��)�r��)�r� �4�dD`���F%H�"�ds�����bT�8L3�(�h&��)�r��(<� ��� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:d`!P̠!��"��G6��9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"����(�̫����)�r���:	@��2� H����������������������A�r��)�6be��3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��e�A3�V����r��)�|�HL3�(�t�d%��2"PȉC"%��2"PȉC"%��2"PȉC"%��2"Pȋq%�8�:P28�� )V��?  �e!M��3�2NS��9NS��9NS�%���3�`�& �0�Qf��i�r��)�*
�8�?�B��$O���@�&Y�H�b��k5�I #,�H&L�@�?�������������������������������������������������������������������������������������������������������������������������������������	$I2d�
%���k�# P(e�d����$I@�P?���(<�9NS���1 �ȫF�`��9�c��9�c��9�c��l 	��/��9h��6�1|�I�r��)�r��)�r� �4�d@��F �<�R�� �J�'	�ze��p�9NS�6@`c>��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�T#�3��9NPygL�*�1�msh�#�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��mP�O h^�/2�e$dr��)�#L�$	F@���"�����������������F���Tq�r��(,و�2#1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q����A3�V�f�@��)�r� ���8(	C"%��2"PȉC"%��2"PȉC"%��2"Pȋq%�8���*�@# A�����7x8 �#&f��)�r��)�r��)��πX,@(�?������U
�TfLə?���X,�9NS�����HR����&L��+ƳY��&L�2��������������������������������������������������������������������������������������������������������������������������������������"I�&000Q(�Mf�X�!�@�,�$����"CC����|�)�r�͘�L�U�p0	��C�1�C�1�C�1�C�1�C6�f��g�	���d��͘�>�$�9NS��9NS��9O�x��Q4�d@��^ Џ�4#�i�ȟ �r��)��σ=3�@�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]
EB>9NS��9L�*�1�msh�#�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh����E�Ṳ���S��9NPH���/AD����������������������*��9NPY�"!<dFbFa?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K����9+/�xW�1r��)�|�HL3�(�t�d%��2"PȉC"%��2"PȉC"%��2"Pȋq t�d*b��=	!T�a� �)
F�h8T 3��9NS��9NS��9A`�X���b�&&%H�!@�P_°���|_
����Car��)�*
�8�?�B�������e�aX�5��d�H```�2aD��"�������������������������������������������������������������������������������������������������������������������������������������$�2c�D�k5��@�P(e�d����$Ha�s*eL�P| �S��9Af�@�&r*Ѹ��!�b�!�b�!�b�!�b�!�b�!�&�	�؂g"��0/�,وdd�Ӕ�9NS��9NS��>�$#8���g1V���)�r��0Y� ��� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:d`!P̠!��h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D�6���x�H��9NS��> `�$	 ^��������������������� ʙS*f��i�r��(,و�2"�f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3	xW�1r��)�|�HL3�(�t�d%��2"PȉC"%��2"PȉC",	ĕa�a"� � p��6e��*�'�<d��)�r��)�r��)�r��i���y��C(eblD!�``` H���B�U `�σ��9A`�Y��~�!K����dɚ�f�Y��I$���,�L�0�"B��������������������������������������������������������������������������������������������������������������������������������������D�	L�2A �$�@F�Y�
�@�������$H�``eL��	A���r��(,و�U�g L�(�1�C�1�C�1�C�1�C�1�C�1�C�0���2;L�U�$^ �l�	�2fi�r��)�r��)�r��A�9NS��9NP,�����H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��*��r��)�d`!P̠!��h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��(W'�4/Q�W# 89NS��	A����~2@�	�����������������BA�4�9NS���1^DU��2��~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����rV_��2"�6b�9NS��> a0�L���2���2"PȉC"%��2"PȊ�d# t�d*q R��q��#A4*��r��)�r��)�r����Tp��q� `�d̙��@�Q(�I�'�� H�T*�P��EA�9NS�Tq���!K����	L�1XV/�f�Y$�2��dɄ	��������������������������������������������������������������������������������������������������������������������������������������ɓ$�I$k5��@�P:��������$H�``eL��	A���r��(,و�EZ L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C73� ��P^�&Ge�dE\f��f�@�#&f���9NS��9NS��9NS��9NPygOM�a��L�f	��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�� ��|r��)�#L鑀�@C2��>M� �m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"����(�̫����)�r�������$O�����������������t	3L�4�9NS�l�	xW3�3	��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>��e�����͘�9NS��*��,_�1*@��'J(dE�8��3 � ����g�8@e��"dd�Ҡ���)�r��)�r��(,3L�4 �3���2�P�2@���H&L�����B�Uњ�σ��9A`�Y��1$O���2̲@�+ƳY��I&L H��"B��������������������������������������������������������������������������������������������������������������������������������������D�&L�H2���V�@�:	�, H����!S*eA�i�9NS���1U��@?�1s�1s�1s�1s�1s�1s�1s�1s�1�`��L���Ȋ��#�͘�>�$�9NS��9NS��9NS��9NP�D��%*c#��g$� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:d`!P̠!��h�#�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m<�x3� 
��Y�r��)P| ����2� H�������������������: f��i�r��(,و�2"�f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3������pY�')�r��(N2��zB��2���'@�B�f0I��I
�3� 'HR4A��2NS��9NS��9NS�F��X,�0�bbbT��R(
�|_d�G����D��T*�h�	A���r����3����)
_����fY V��XV/�$��H$&L H���������������������������������������������������������������������������������������������������������������������������������������$�2fY�H�b��k5���H$�����#*eL�,9NS���P&*�Xp���C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�3s1� 	���dv �ȫC0�����l���r��)�r��)�r��)�r��M��$FK�/ �L�f	��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �WB��P���S��9NS#
��exB�����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� ����m2��ʹ�Y�r��(J> H2@�	�����������������
 @�3LӔ�9NQ�b�2"�f!�f����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3	xW�1r��)�r��f�g1Vq��M��d��l��UDM��2����)�r��)�r��(<�3���3�0?������؛b)
B�$�'������B�UњT 3��9A`�Y���!K����dɊ±|k5��$��H$&L H��������������������������������������������������������������������������������������������������������������������������������������$�2��D�k5��f�A �����D���H @�,9NS���1UJ��	����9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c�� ��P^�&Ge�dE\f��p� &�ə�)�r��)�r��)�r���&2c,	�HR�W��`��e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�T#�3��9NPygL�*�1�msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&�G6��&�>� �����)�r���$	 ^��������������������� �i�f��)�r��8f��s1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��Q�K�Ȋ�,و��9NS��	A��	��<H�M
��r��)�r��)�r��)�!0L
鑌�bbbfLə
�Y��2�����$U
�T3FhP| �S��A�~?�!HR'����d�A��k5��d�H```�2dɓ��������������������������������������������������������������������������������������������������������������������������������������	$I�e�
%���k5��d�A�������k `� �X,�9NS�g�@���`�?�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���(��L��|���pp��P��4'Ô�9NS��9NS��9FH&��a4)�A�%*c>���9 ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��*��r��)�d`!P̠!��h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D�6��� d�H��9NS��> `�$	 ^��������������������� �i�f��)�r��8f��s1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q����A3�V�f�@��)�r��)�r��)�r��)�r��)��σ$G̐�g���e��Gdv��P(``` H�������$H�B�f�� �|�)�������)
_����fY V/��X�/�%��H$&L H��"B�������������������������������������������������������������������������������������������������������������������������������������� H�dɌI #Y��k5���/����	k5���3�,9NS���1U��@?�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1��r�^g�xWٕ�1|�I�r��)�r��)�r���:2A4��LGB�	 JT�|3�29�&rds0L䀲�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�T#�3��9NS���B�!�@C&�G6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��mP�O h^��2e$dr��)��πH���/AD�����������������5��f&&&H��#��9NSdd���2"�f!�fHϸ���\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\9�`�{2�hN�)�r��)�r��)�r��)�r��(<���a0L  	���0g�2fL�@�P(�J$ɓ���������"A�x3FhJ>S��A�?��!HR����D�fY V��Y��I$���A �2aD��������������������������������������������������������������������������������������������������������������������������������������@�$ɓ$�I$+
��|_
ĂA�������k `� �X,�9NS�g�@�W���2�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C73� ��P���^DU�����ə�)�r��)�r��)�r���:2A4��C"U� 4φy�G3�H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�O��G�g)�r���4ΙT3(c��"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m<�x3� ɔ���r��)�	@��2��������������������������$r��)�l��� �ȫFrV_�����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������J��"�D���r��)�r��)�r��)�r��)P| ��4� �0�?���2���6 �P(�I&O��������$U
�T3Fh<�3�)�r��`����)
B�����ɓ����k5�I !���dɄ	$O�������������������������������������������������������������������������������������������������������������������������������������D�	L�2A �$�@B��_�f�A �����D��f�X,r��)�F��+�bbds01s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13�������^ NS��9NS��9NS��9NPygFH&��a4e�"2X�,�9���3��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�O��G�g)�r��)���@C2��>M� �msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D�6��� d�H��9NS��> `�$	 ^�������������������+
���">d�S��9HМ3�Ȋ���Q�O�������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������C(�&rV_�129�	���3�x>�$�9NS��9NS��9NS����t��$8㘘���2fE�A��k&L����������$U
�T3FhP| �S��A�?��C�	���̳,�+
���k$��FY �L�0�"������������������������������������������������������������������������������������������������������������������������������������� H��"I�,�I��k5���, H����k5��LLA`�Y�r��)�`�� &b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���|��0/�2fi�r��)�r��)�r��)�r��$A�0��2����>����*��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:d`!P̠!� h^�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD͢'�4/}�2�29NS��	A��$	F@���"�����������������±|bbbd���9NS��#Bp�L�U�1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\f!�f1�0���P����g"�"���f NS��9NS��9NS��9NS4�3Fh�?���(e�;#�D�!H�I	����������$U
�T3FhP| �S����g���0�?����Y�H�b��k5�@@#,�H2̲@@�?��������������������������������������������������������������������������������������������������������������������������������������"B�$�H2�$�|_
ƳY��H2����(�J%�_��f��i�r��)�`�������1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��$hN�)�r��)�r��)�r��)�r��(g�0��2%\��Xφy��fJ����� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:d`!P̠!��h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D����"�*�RF@g)�r��(<�� H��$O�����������������X�/�LLL�2G)�r��hN�	���+�$<������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFa3��������	�"�1 ��+�	�2fi�r��)�r��)�r��)��0�@�"te�@�PQ(�I�'������������	*�P��4%�)�r��`����b����dɊ±|k5��  ���2d���D�������������������������������������������������������������������������������������������������������������������������������������$H@�$�A�I$����V�b��H2������������4�9NS��#Bp�ٕ L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C73�9�`	��\��g�@��9NS��*�J|��P_���r��)�r��)�r����3��>g�8e�"2X�,g�<�� dB�@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]
EB>9NS����t�h�  ���&�G6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh��m2��ʹ����r��)P| � H2@�	������������������k5���#�H�9NS��34A3�V�t$������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.���H��e�s���>J�V���6�1l����σ��9NS��9NS��9NPX,��y�blA�t$	������������$H�B�f��"����)��� H1����2d�aX�5��d��$	�&$H@�?�������������������������������������������������������������������������������������������������������������������������������������	$I2d̳,�000+
��|_
ĂA�����$/��/�4�3NS��9M��3A��eM�2�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��)�#K�� ��  '���T����)�r��)�r��(l���g,	��xc>��"��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�O��G�g)�r���d� �S8#� g�ɴD͢ �msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴDB�<�x2��ʹ����r��)P| � H2@�	������������������k5���#�H�9NS��34��`�䬿���q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFa3����&��
��@���	�0�> g)�r��)�r��)�r��)�|�H �	��2�(
2̲@@�?�������������	*�P��4�> g)�r����b��C����	e�d�XV/�f�Y$�2��dɄ	��������������������������������������������������������������������������������������������������������������������������������������D�	e�d�I$+
���k'����@@"�/��3L�4�9NS��34f�����`b����C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nc=2B��Hx�l��� ��*���
��r��)�r��)�r��$A�̪��`b�xc>��"��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r���:	3�< z|�DA�"|�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh��m3� 
񔑐�r��(J> H2@�	������������������/�c?��0L�)�r�#&f�R�9�����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��2��9�e�dvUJ��H��,وdd�Ӕ�9NS��9NS��9NS��9NS�Ca_��_ƳY���������������2d�P�C4f���:r��(l�,P(�����Y�H(�J&�Y��I&L�2�������������������������������������������������������������������������������������������������������������������������������������$I2d̳,�000+
��+�D����H2�P�2D|��)�r�#&f��0/�^g��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�AW71#Bp�9NS��*���������`N2�0�L� ��A6fdf
�`T�@J|�A�9NS��9NS��9NP�|2�* e�����y%� 2!] ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�O��G�g)�r���d� �S8#� g�ɴD͢'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DA�"xB�ey�s)# 3��9NPygA H2@�	������������������Q(���2�`�&9NS��6FL�*�Xs1�0������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\~>������q��\f!�f]	!�3��D'��W�����>*�)�r��)�r��)�r��)�r��)�r���9�6&ę2���������������B�Uњ�σ��9A`�YbŊ�@�?����2b��_�f�I$000L�0�"x@�?�������������������������������������������������������������������������������������������������������������������������������������	L�2A �$�@E�D�k5����I$��P�FH��#��9NSdd��p��P<�ϑ�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nc) #/5���@@ơp�&�̌�P
��#O��T 3��9NS��9NS��	A���*��X���Ы@�71VX���� ,�e�,@Yb�X���� ,�e�, �WB��P���S��9A�i����=>M� �m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"�\� мD^e\�H��9NS��> `�$	 ^�������������������Q(�FP�A0L�)�r�#&f�R�9�����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3�!��	��xW�`_�Y�'�<d��)�r��)�r��)�r��q)�c&)�c&2A4r��)�r���:~?��@@�?���������������B�UњT 3��9A�i�,X�@�P'����&L�Q(�±|I$���,�L�0�"B���������������������������������������������������������������������������������������������������������������������������������������	L�2A �$�@B��_�f�����"�������C(&	�c��9NSdd�јF�����1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r���P_�8,�� ���j5���@@ơp�&�̀�b*ʠ%> ����9NS��9NS����tٕQP�G�e��g�: �W@�
�e�,@Yb�X���� ,�e�,@Y` dB�� ��|r��)�#L�$�3���"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m>M�&Q�W2�29NS����t�~? ^�������������������Q(�FP�A0L�)�r�#&f�R�9�����}.?K��������}.?K��������}.?K��������}.?K��������}.?K��������}.3�3	��Q�L䬿�	��!<dDd3����	�0�����9NS��9NS��9BPy�*�3ќ2��,g����=�͑�r��)�~?��@�?��������������� B���@�4Μ�)��"ŋ
��"���2d�aX�5��d�H�$	�&$O��������������������������������������������������������������������������������������������������������������������������������������	L�2A ��b��k5�I /�������#�H�9NS��34f����>G1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�?�
���ϊ�1�r��)P| �8,�� ���j5���@@Ơ cP��!Ђl���#8X%> ���)�r��)�r��(l��UM�aV/$��a D+�� ,�e�,@Yb�X���� ,� 2!]
EB>9NS����t
gx@��6��9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h�#�DO�h��� W�����S��9NS���d�z'�����������������D�QC(er�FNS��9O�x�*��"�C���\~>������q��\~>������q��\~>������q��\~>������q��\~>����bFa3�3�!��	�؂g"�"���f M��3J��r��)�r��)�r���4΄���S��L��f�*^�U�ye����lD`A �6eTT9NS����t�?�
 �"��������������	*�P��4�> g)�r��`�ŋ
���ɓ&+
��+ĒH```�2dɓ��������������������������������������������������������������������������������������������������������������������������������������	$H@�&Y�H(�J&�Y�``` H����I$�����L�)�r���<d�"���dv9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c�� ��PU��F|T	�S��9J��)�`le e�@Ơ cP1��j5���@@Ơ cQ����&�̃
s`
pX��W*��r��)�r��)�r��qlʨ�zn3 �/䗐l  ȅt���� ,�e�,@Yb�X ��?�"���)�r���:	3�< z|�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴDB�<�x2��ʹ�Y�r��)P| ����2� H�������������������De��Uʹ9NS��>�$�����I'��q��\~>������q��\~>������q��\~>������q��\~>������q��Q�L�2�� ��P"�D+�b8W�Y�'�<d��)�r��)�r��)�r��M��=�LGB�! �nb�6"0�!%��VR+)?��X�䗐l$|�Fq�r��)P| ����@�P'��������������@�"�U
��3@�Py�r��(<�3��(
����&L�Q(��f�I$e�	ɓ'�	�������������������������������������������������������������������������������������������������������������������������������������@�$ɓ2̲@����+ƳY��I	�������L�)�r���<d�"���dv9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c�� ��PU��F|T	�S��9J��)�`le e�@Ơ cP1��j5���@@Ơ cP��4�Hx�l��0�6 ���d ���9NS��9NS��9BPy�lʨ��dU�GB����X@Yb�X���� ,� 2!]
EB>9NS����t
g	���msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&�G6��&�? ����)�r�����# d�@�?�����������������%��C(��r2r��)�|�IU*�3��I'��q��\~>������q��\~>������q��\~>������q��\~>��e�s���쪕`�a�'���*��r��)�r��)�r��(l��UM�`�"��:hds0L�� ��e'��YI����VR$�V�/ �H�����9NS��?�
 �"��������������	@�3��3@���r��(l�,P(�����D�±|k5��$��H$fY  H���������������������������������������������������������������������������������������������������������������������������������������D�	Y$��b��k5�	�����#�Cc��9NS�2L�xb�2;�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A��6/0W @Ơ cP1��j5���@@Ơ cP��4��X&�8^���
� Fq������T��9NS��9NS���͐�	����dU�^Iy� �WH,@Yb�X ��?�"���)�r���:	3�< z|�DA+���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m>M�&}�# 89NS��9A H2@�	������������������Q(��8G0��)�r���<d�ss]	!��}.?K��������}.?K��������}.?K��������C(�&rV_�a �L�Bxȅx�@ �
�IDhN�A�9NS��9NS��9NS�F��P���a4e�"2X�,�f*�`� #����O�Z�=*�5�YI����U�j3ҭQ���X�䗐l$|�Fq�r��(J>���@�P����������������B�Uњ�σ��9A`�YbŊ�����ɓ�b�V��I$000L�0�"�������������������������������������������������������������������������������������������������������������������������������������D�	L�2A �$�@E�D�k5�I  �"����e��#����9NS�2L�x`<�ϑ�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 2�d��R F^j5���@@Ơ cP1��j5�`N3A�81��j5����L����8Xg͐�T 3��9NS��9NS��	A���	�����T��^A��"� dB�lD` dB�� ��|r��)�#L�$�����mP�O�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��(W'ɴDϸ #&RF@g)�r��A�� H��$O�����������������D�G� �@��)�r� �U��Et$������}.?K��������}.?K��������C(�&bFa�2�2;L�U�$^ �l�	�2fi�r��)�r��)�r���4΀�f�S��L�HU�V�	
� ,��!%��VR+)?�����O�e'��YI����VR*�5��!%��^Iy�G��g�)�r�����P(	�������������� H�B!�њT 3��9A�i�,X��P('����&LV��Y��I$��	�&$H@�!D��������������������������������������������������������������������������������������������������������������������������������������"B�$�H2�$�D�Q5��d�H H����e�d�8G����> g)�r����6/`#��C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nb�3rj5���@@Ơ cP1��j5�`N3A�3����j5�`Njў�!_A�9�8,�a(|��9NS��9NS��9BPy�)�c&FFh&�?�$t*�< �� ��2����9NS�S���
gx@��6��9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h�#�DO h^��2e$dr��)��πH���/AD�����������������(�J$p��
D	�r��)�%\��WFA0?K��������}.?K�������3�"g%e� L�(	�"ٕ¼ ��� �r��)�r��)�r��(<�3�1�F��=�,	��x`71Vd��X+)?�����O�e'��YI����VR+)?�����O�Z�=	!�g�y%�	3ќr��)�T 3���a&�D��������������$U
�T3FhJ>S���͑bŊ�@�?����2b��_�f�I$e�d�dɄ	��������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$�D�Q5��d�H H����L�28G����9NS��> e��W��2;�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A�/�L�e e�@Ơ cP1��j5���@@Ơ cP��f�p cP1��j5�h0'���D/Fzd�}��/�L�	@2����)�r��)�r��(J>8Ld���Ч��R�FFh&��f��9NS�F��H)�� 3���"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� �m<�x3� ɔ���r��)�	@��2������������������(�J$p��
D	�r��)P| ��g�]	!��}.?K��������}.3�3����^�&Gb	���d���p��#&f��)�r��)�r��)�r����S��L��f
�*؁#�V���fJ�� ��e'��V���J�O�e'��YI����VR+)?�����O�e'�Q��h��$�ɟE䗐l$|�Fq�r��(<�3��$	 ^��'�������������� H�T*�P��A(<�9NS��,X�P(���L�2�D�k5��$��H$&L H��"������������������������������������������������������������������������������������������������������������������������������������$ H��"I�,�IJ%Y��I ������ɓ3&d̀P
 J��r��)P| �����dvnf9@s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�?�
���ϊ�1�r��)P| �8,�� ���j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'`�d#,�@��	 ���0�>
��r��)�r��)�r��(<��ٕQP3�Ӕ�9NS�F��H)�&g�ɴD͢'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DA�"|�DL��2e$dr��)�T 0H���/AD�����������������(�J$p��
D	�r��)P| �x�@ ��r���\~>�F}�$L䬿�bds0BxȈ�g��z+�,و����)�r��)�r��)��ρP���a4dJ� � f��� t�<�A	,U����YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�Q����3輒������9NS����t�# d�@�?���������������B�UњT 3��9A�i�21��t�P(���L�2�D�k5��$��H$&L H��������������������������������������������������������������������������������������������������������������������������������������$ H�,�$I "�D�k5��  @�?����2fd̙� �S��9J��_�E/`#�s1���9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c�� ��PU��F|T	�S��9J��)�`le e�@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N3A�8�8^�	 �)̀)�`l	@3�/�)�r��)�r��)�r��)�r��(<�3��S8L�O�h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D���ϸ #&RF@g)�r��(<�� H��$O�����������������D�G� �@��)�r��W����&�2��9�e�dv �ȫC0�����l���r��)�r��)�r��)��#fUE@8� ����Z���*�`� #����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�Q����3輒��&3NS��9NPH���/Dɓ��������������$H�B�f�� �|�)��"ŋ
 �"���2d�aX�����I&L�2�������������������������������������������������������������������������������������������������������������������������������������$I2d̳,�I$��%���k$��AD����dɕ"�T�0��t�9NR�����_����s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13���������)�r��S����@����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j���f�q�	�X&�8^����W3M��ɟ�a(|��9NS��9NS��9NS��9NS�q�*�
���#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD͢ �m<�x2��ʹ����r��(J> H2@�	�������������������2f@(')�r��(<�2E��X�0��2�,��&x3��Q�aP| �S��9NS��9NS����td�h<���� �a��0@q͂��C�Ϣ���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR*�5�V���J�O�|3�	�LӔ�9NR���@�$d�z'��������������@�&�؛<�Py�r��(l�,P(�����ɓ(�J&�Y��I&L H�$O�������������������������������������������������������������������������������������������������������������������������������������D�&L```�IJ%Y��Q(�I�'���ɓ&fLə �0F�Ӕ�9J��gT$��2;�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A��62�2� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơ�	�h0'���f�
f2�0�D	 8_�|�3�% ς���)�r��)�r��)�r��(� F|0�Ȭ�&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��msh�#�DO�h��E�Ṳ���S��9J��	@��2� H������������������H�  �S��9NPY�#8W�Y�&�ə�A�9NS��9NS��9NS�%��&2`p2AO�	y%�	y���6"1YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��V���J�O�|3�	�LӔ�9NP�|@�$d�z'��������������6&�؎8�(<�9NS�6FF20��
 �"���2d�aX�����Q(�d�A2d��'��������������������������������������������������������������������������������������������������������������������������������������"B�$�H2�$��+ƳY��Q(�	���ɓ&T��R �0�9NS��> c8W��2;73�9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��\��g�@��9NS��*�~2g�) #/5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���C4��`Nj`�d"��3Epl�H 2di{>
��r��)�r��)�r��)�#L�S��1 3�Xq��G6��9�D͢ �msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DA�"xB�ey�r0����9NPygA H2@�	�����������������```�"��`�r��)�r�����9NS��9NS��9NS�d�h<�����! �|3�2�� �&}��ʴFzU�j3Ҳ��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�Z�=+)?��� t&3NS��9NS���d�z&L����������������"M��6#�8J>S���͑bŊ�@�?����2���_�f�I$e�	ɓ'��������������������������������������������������������������������������������������������������������������������������������������@�$�A�I$��%���k(�J$ɓ����ɓ*EH��x#L��r��)�P�������r��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR���pX��+� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'���e�a��>Dd��~2g�&F���/�A�9NS��9NS��9NPygH����? �� 3���"��G6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��9�D�6���x�H��9NS��� H��$O�����������������Y��G��C�)�r��)�r��)�r��)�r����S��L��f
�*؁#�V���fJ�� ��e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3ҭQ������g�:��)�r��A�� H��$O��������������lM��q�Py�r��(l�,P(�����ɓ�b��k5�I #,�H2̲@@�?��������������������������������������������������������������������������������������������������������������������������������������"B�$�H2�$�|_
ƳY�V���"���@� �C<��<�9NS��> fpUBJ����!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�AW71�P&9NS��*�����������@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N3A�8��!/0W$d���  d���A~9NS��9NS��9NS�S����L��ɳ3� 
�=<�xsh�"�p"|�DO�h�#�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� ������E�Ṳ���S��9J��~?���/AD����������������L�3Y��P(ə3'����3LӔ�9NS��9NS��9NS�F�ђ	��>g�8,X�,g�<��(�	!�g�V���J�FzVR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�Q������g�:��)�r��(<�� H��$O��������������lM��q�Py�r��(J>,(
?���&L��+°�_I #,�$fY  H�$O������������������������������������������������������������������������������������������������������������������������������������� H�A �$�@E�D�k5�±|$O���$U
�T��y�r��)�gT$��2�,s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13���������)�r�A~�6/0W @Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơ�	���@@ơ�	�Be e�d��~2g�4�*�A�9NS��9NS��9NPygE8�>
��Ɂ���3? �� 3�����"�\�(W'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&�E
�D�6��D^e\�H��9NS�%������$O��������������ɓ&I$��@�Q�2��}>���� ��4�9NS��9NS��9NS��> `0Y���H)�A#�V��G3�M���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�h�����g�<�ИD�9NS��9GsblM�2d��������������� d��T 3��9@`�dX�b�@�����2d�%��+ĒH�$	�&$H@�?��������������������������������������������������������������������������������������������������������������������������������������"I�&H$d�H�Q(��f��D�L�?���$H�B� M��9NS��¼ ���af�c�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13�������8f�)�r��S��ؼ�\����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��2�0�D	!�* A�T��9NS��9NS��9NPygE8�>����? �� 3���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD����"�*�RF@g)�r��)��~2@�	�������������� H��D�b�"� ��p�&	�`�X<�3�)�r��)�r��)�#L�l������1c<� 
���@F$�V
�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��V���J�FzVR3�@�L"f��)�r��q�6&�ؓ&O��������������6&�؎8�(<�9NS�6E�(
D�����"EaX�5��d�H�$	�&$O��������������������������������������������������������������������������������������������������������������������������������������	L�2A �$�@E�|+�f�XV/��'�����B� M��> g)�r��8/c,eY���!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR����&2�2� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơٙ���A�9NS��9NS��9NS��9A�i��$�# 8?�_���G� �O h^�h��msh��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h����E�Ṳ���S��9J��	@��2� H����������������F�؛�2�Q���4��$T 3��9NS��9NS��9A�i���H)�A#�V���fJ�� �� ��*�V���J�FzU�j3Ҳ��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3В&}�� t&3NS��9BPy�+�F21�6&ę2���������������6&�q���t�9NPX,X�a@�Q����2d�aX�5��d�H�$�,�$H@�?�������������������������������������������������������������������������������������������������������������������������������������	��$�I$Q(�Mf�X�+�ɓ����D���  �<�3�)�r��8/c,eXg�@�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR���pXHx1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cQ����1� ����)�r��)�r��)�r��)�r�q�|���/�~^L�O h^�"����"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴDB�<�x2��ʹ����r��(<�3��$	 ^��������������&L�D�Q(
d̙�H�0���X,�9NS��9NS��9NS��	A��L"f��*^�g�:e�A$>L�+)?�h���@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�h�����g�<��8�#��9NP�|8�vG`�L�?��������������؛b8���9NP,�,XP(���L�1XV/�aX�$�@FY �e�d��"x@�?������������������������������������������������������������������������������������������������������������������������������������ H��"B�$�I$Q(�Mf�X�+�ɓ����؛b8���9NS�'��e��7 ��1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nc) #/5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j�� �J|�)�r��)�r��)�r��)�r��)�)�I�e$d��x@A3=<�xsh�#�DA�"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��mP�O�h��E�Ṳ���S��9J��	@��2� H������������D�I  P(d�z>�O�TʙQ�3@��4���t�9NS��9NS��9NS��9NSfUEB�xc`� #����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�Q��h������f*�8�#��9NP�|
鑌�lM��&L���������������lM��qʃ�r��(l�,P(�����D�±|k5��$��H$&L H���������������������������������������������������������������������������������������������������������������������������������������ɓ$�I$+
���k5��dɓ����D�blL�da]	A���r��(��D'����r��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR���pXHx1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���C4��`N"��*���S��9NP�|
�|)�c&*�J>S��9NS��9NS�S����H�
g~^L�O h^�"��G6��&�G6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD�6��&�(�̫����)�r�����~? ^�������������&LV/�����C<111q�`�&��`�4Μ�)�r��)�r��)�r��)�r��p2F|3�+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��V���J�O��*��<���:r��(J>sblM�2d��������������� d��#L��r���X,�b��C����,�$
±|k5��$����2dɓ'��������������������������������������������������������������������������������������������������������������������������������������D�	H$d�H�Q(��f�XV/��'�����6&���FД|�)�r�͘�	�"73�9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��\��g�@��9NS��> b��R F^j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�f�qp��P��8r��)�r�2�*?�%��2�O�L"f��|#L��r��)�r��)�#L�'�� F|
g~^#� g��4/ɴD�6��9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M�'ɴD����"�*�RF@g)�r��)��~2@�	���������L�1���t	@�����?��h�2D|��`���9NS��9NS��*�P| ʃ�r��)�r��)��p3aYI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���ʴFzC�Ϡ71V�<��)�r��q�6&�ؓ&O��������������6&�؎8�A�9NS�F��ŋ
��"���2d�aX�5��d�H�$	�&$H@�!D��������������������������������������������������������������������������������������������������������������������������������������"B�&L��e�	$�D�Q5��f�Y��2��� H�blM����+�A�9NS���1"�Dnf9@s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�?�
����a�r��)P| ��?�Hx1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơ�	�A��3@0� ��r��(<�3�p2Dt*�< ����� �����23A4T#�0ygNS��9NS��9NS�S����H�
g g�8  ��� м9�D�6��&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h��m>M� ����m3� 
񔑐�r��)P| ����2� H��������� H��D�b�"� ��,!�0�A�r��)�r��)�r��)P| ς��24��pX�����8r��)�r����0φy�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR*�5�YI���U�p2G)�r���4Ζ,X؛bL�?��������������D�blGp�|�)��"ŋ
���ɓ&+
��+ĒH�$	�&$O��������������������������������������������������������������������������������������������������������������������������������������	$I�e�	$�D�QAАk5�ɓ'�����2�� �|�)�r�͘�	�"73�9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��\��g�@��9NS��> b��R F^j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�f�qp��P��8r��)�r�����H,@Yc#��g nb�#�V��O�̐�	��<�3�)�r��)�r��)�#L� F|
g g�8  ���dVA�"�\�&���"|�DO�h��m>M�'ɴD�6��&���"|�DO�h�"�p"xB�ey�s)# 3��9NP�|@�$d�z'��������@�Q�6&��}>����<̑2EA�9NS��9NS��9NS��> c>l��, Fq��l����!$|I�  �*��r��)�zn3 U�+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��V���BH|���f*�8�#��9NS� M����	�'���������������blGp�|�)���,P(�����ɓ(�J"��_I !���dɄ	$O�������������������������������������������������������������������������������������������������������������������������������������D�	$I�e�	$�D�Q5��f�Y��2���� ^����P| �S��9Af�@���sp0	��C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A��6/0W @Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���B �z��	O�p�9NS�� ��� t���� ,�e��f	�������Z�?� p2B�&2a(<�9NS��9NS��9NPygL���� �p }�	��E`�6��(W ���"�p"|�DO�h��m>M�'ɴD�6��&���"|�DO h^�/2�F pr��)�T 0H���/AD�������dɔJ%�@�T��R/��/�ŋr�FA`�Y�r��)�r��)�r��A�	O�pɑ��3�W3M��f
���yM�M�hUJ� �32	@3��9NS���f�� t���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�Z�=+)?�����H�9NS����<U
�TL�?��������������؛b8ㄠ���9NPygK,P(�����ɓ(�J&�Y��d�A2d�����������������������������������������������������������������������������������������������������������������������������������������"B�2̲A$�(�J �:f�Y�e�?���@�"�@��?�����9NS�l�	xW7 ��1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 2�d���f
��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�D/F�d� ��S��9BPy��3�@�e�,@Yb�X���� D+�t*�<U�V�̐�	��l�S��9NS��9NS�F�� ��$� �#�C2��Ȭ� м(W ����m>M�'ɴD�6��&���"|�DO�h����E�U���S��9J��	@��2� H������ H����t	@��8G�2�T �34�3A�i�9NS��9NS��9NR�����>
�����"	�3#4S0��L�A��F�z4sѠ	U*�x��2di{9NS��9OM�a��J�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3Ҳ����� �d�S��9NP<ʑR*Dɓ��������������͉�6#�8J>S���͑bŊ�@�?����2b��_�f�He�	Y�H'���������������������������������������������������������������������������������������������������������������������������������������&L��e�	$�D�Q5��f�Y��2������I����~��t�9NS�l�	xW7 ��1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nc) #/5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��3A�8�8^��� )��)�r��`c>��X���� ,�e�,@Yb��9p3a
�dU�zn38Ld�Py�r��)�r��)�r���:#L�L_�R��`�`!�@C м м&�G6��&���"|�DO�h��mP�O h^�/2�e$dr��)��σ���d�z'����ɓ&I �C�"�T�LLK,!�0���a(<�9NS��9NS��9NR���A~��~2g�8_�|�@�ʜ���*�S7E4sѣ���h�G=n �ix��#>F')�r���4Ξ���@q��O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3Ҳ����� �d��i�9NS����<�"�L�?��������������؛b8ㄠ���9NP,�,X�P(���L�1XV/�f�Y$&L�@�< H���������������������������������������������������������������������������������������������������������������������������������������&L� �e�I "����t$��H$����$H�P(?����4Μ�)�r�͘�/"*�	����9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�f�c� ?�
���ϊ�1�r��)�T�Nc) #/5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��3A�8�8^��� )��)�r����,g�<���X���� ,�e�,@Yc(� ,�e���X^Iy�L�x=7��&2`�4Μ�)�r��)�r��(l�3㈄�0�0̠!�2+ �ɴD�6��&���"|�DO�h�"�p"xB�ey�s)# 3��9NP�|@�$d�z'����	L�3Y��d�z>�O����f��#$G̐J>S��9NS��9NS��> eA�	O�pg � �bg�HWњ)�P8
7E4sѣ���h�G=9���F�z4�A��3r2F|�NS��9NS�q�g�<�Ҳ��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�nb�=7�)�r��(��H�"d����������������@����> g)�r��f���Fҁ@�$O���$�Q(��f�He�	ɓ$ H���������������������������������������������������������������������������������������������������������������������������������������$�2fY�H�b�BA��k$����$H�P(?���A�9NS���1 �ȫ@	����9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c�� ��PU��F|T	�S��9J��)�`le e�@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'ѳ  %>Ô�9NR�������H,e�D� ,�e�,@Yb�X���� ,�e��
�y%�2����f2�*����9NS��9NS��9A�i�@ϙT �3\�UȬ�9�D͢ �msh�#�DO h^�/2�e$dr��)�#L�$	F@���"��L�2�D�P(
�R*F&&%� �@��`���9NS��9NS��9J��|��e�ɟ��~	��3rT�d��	U*��G=9���F�z4sѣ���h�G=9��qSK�����19NS��9@�d��g�:C�Ϣ���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR*�5�YI����T��Ô�9NS� M��g�ɓ��������������͉�6#�8J>S����t�b��C����,�$
±|+
��$�2��dɄ	��������������������������������������������������������������������������������������������������������������������������������������D�	e�d�I$+
��(
AА001�����P(?���(<�9NS���1^DU�?�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13���������)�r��S����@����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N"�f2@ J|�)�r���4Ι����H,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]/$��a�T� e���U `�dr��)�r��)�r���4Εs$F�AL�0�rTS"�
|�DA�"����(�̫�I��)�r���# d�@�?��@�Q�2��8eL����<��$r��)�r��)�r��)�T 1�6B�� #8�A6fdf�
fl%T�����z4sѣ���h�G=9���F�z4sѣ���h�M�M/0W!8NS��9NP�D�/$��a	!�g�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O��fJ���f��:r��)���yR*EH�2���������������6&�؎8�A�9NS�6E�(
D����dɔJ%Y��I$���A �2�ɓ���������������������������������������������������������������������������������������������������������������������������������������"I�&H$d�H�/�`t	 �:	�/����	bʙS*�σ��9NPY�"	��� ��P9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��\��g�@��9NS��> b��R F^j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�f�qp�1� S�9NS��	A��Xφy�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�䗐l tʗ��q�lʨ��#��9NS��9NS����t��"4q�fD^e\S"�
|�DE2+ � g�8 ��9NS��	A��bŌ��/AD�L�2�D�b�g��_��X�a!�0,9NS��9NS��9NS��> g�P_��^��?�s4�e e�NFK�n �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)��f
�'���r��(<�3�p2E䗐l%e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����̕A��9NS��*���H�"d�����������������؛���)���,P(�����ɓ(�J&�Y��I&L H�$O�������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�aX�AАk5��?����!H� �X,�9NS�g�@�A3�V�?�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13���������)�r��S����@����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N"��* @J|�)�r��)���� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+� ȅt�������e���U `�dr��)�r��)�r���4Ίq�|"��#�(�̫��x
g�d�)�r��(��d̙��D�e�	�Y���}>�O����fH��"����)�r��)�r��)�T 0��p<��bg�HWњ)�P8
7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4�@��p<��)�r��df�iy%�I�>��O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR/32U��0F�Ӕ�9BPy���x!�	�'��������������� ^�p�|�)�#L�bŊ�@�?����2b��_�f�I$e�d�dɄ	$O������������������������������������������������������������������������������������������������������������������������������������� H�dɒ	Y$��b�
��H�����k5���2��4�9NS��6FL��1 �<�ϑ�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A��62�2� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơp�1� S�9NS��	A������ t���P�$@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yc`� #��*� dB�g�<�Ҭ28�6eTT�͑�r��)�r��)�r���:��� �,� �,S����9NS��9L�4�?���D2�˦d̙�ŋ P
 EAPg�)�r��)�r��)�T 3�/�0�/�L��O�HyS���%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSDA��3�b�r��)�r���	�䗐l%e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����̕A����t�9NS���T��2d���������������blM���σ��9@`�dX�b�@�$O���&L��+ƳY��Id�A2d�����������������������������������������������������������������������������������������������������������������������������������������"B�$��������t$��H�����$P�@x�����9NR����p����p���C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�₮nb3�Lr��)�T 1Nc) #/5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��jѳ  %>Ô�9NS��G�g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�y%�	V ��=�0Y�9NS��9NS��9NS��9NS��9NS��2D|�њ3Fh�#�HF�Ӕ�9NS��9NS��9J��3��A�2�g�&�̌�L2�pn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4D/C8X�9NS��##4K�/ �J�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���*��q�r��)�r�`fLə2����������������؛b8���9NP,�@�$P(�����ɓ�b�V��I$000L�2d����������������������������������������������������������������������������������������������������������������������������������������$�2fY�H/��XB@:�����������E�_���1�r��)�%��W��EZ���g�@�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�AW71�P&9NS��>
��_�����\����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���ٌ� � ��r��(J> 2��|3� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y���/$��a*�#�``cfUE@,��)�r��)�r��)�r��)�r��)�r��)�r��)�r��)�r���8d���_���S� ��\��`Nn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�8^�p��r��)�FFh&��^A����3謤�VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��3%Pzn3�i�9NS�� �0̙�2L�?��������������D��T*��<��t�9NQPT����R�/���ɓ&Q(�Mf�Y$�2��dɄ	��������������������������������������������������������������������������������������������������������������������������������������� H��"I�,```V��t	 �:?����ɓ2@����4�3NS��9J��6bf���Ȋ�^gɸ��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�AW71�P&9NS��*�~2g��3rj5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�f�qp�1� S�9NS��9L�ppφy��2��"�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "�>��3�� e������,���:r��)�r��)�r��)�r��)�r��)�r��)�r��A�	O�pg �tf
�`A6fde�a����qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�p��c��9NPygBa4��Z���3謤�VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��3%Pg���)�r��(�fd̙�,�H��������������I ��eїD0��A�9NS�&	�b�/��5������	+
���k$�@FY �e�d��"������������������������������������������������������������������������������������������������������������������������������������� H��"I�,```�/�`t	 �P(�H2������Q(��2f@09NS��9NSdd��Y�#0��^DU����3����r��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR���pXHx1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�8^��� )��)�r�����G�g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����/32U|3�,g��`H��2�* �f��9NS��9NS��9NS��9NS��9NS��9J��|��b���R F^T�d��	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4D/C8X�9NS��	�L�:hVR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI���`�ɞ���:r��)P| �02!�F]2���������������&L�@�P2�Tʂ�`���9A�i�,X��6&��$?���&L��+°�_I !���dɄ	��������������������������������������������������������������������������������������������������������������������������������������D�	H$d�H�/�`t	 �P(�I����D�Q#�p� P
 NS��9NS��9M��3Bp8^���eK�Ȋ�^gɸ��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�AW71�P&9NS��*�����������@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���f
�� ��r��(J> 2��|3� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅtφy���2�,	��D���4%�)�r��)�r��)�r��)�r��)P| �S��2�g�&�̌�L2�pn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G="��Ӕ�9NS�����#�V��$>L�+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����``ygNS����t �32fL�2d�������������$�2b��)�� ��9NS�2@�<#�p��f�����2d�aX�5��d�H```�2aD�	$O�������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$�|_
��:@�Q$������&LP(���PT�)�r��)�r��)�l���3�x�`_��2"�^�&Gf�`��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��\��g�@��9NS��> b��R F^j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��"��* @J|�)�r��)���� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅtφy���2�,	��D���4%�)�r��)�r��)�r��)�T�&F���d��p��x�����*�S�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSDA��3�e�S��9NR>g�8��Z�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR2��!���J>S��9@03&d̓&O�������������
B��*�P� `� ���:r��(<���<��8��  H�����2d�aX�5��d�H�2�ɓ'���������������������������������������������������������������������������������������������������������������������������������������$�2��|+��H�D�H����k5��P�E\�����9NS��9NS��9NS��34'��W���Ȋ�{ ����Lb�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�&ss�c��9NR���pXHx1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�8^��� )��)�r�����G�g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���T ��X�,2��#�z3�`�dr��)�r��)�r��%>�PU0T	�3" �z
F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�і	�B)�`lr��)�r��&i
�	!�g�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�P�$���t�9NS� �3"te�,�H�����������ɓ&+��@�P*EH����8�H��"����)�������P(&L������&L�Q(��f�I$e�	ɓ$ H���������������������������������������������������������������������������������������������������������������������������������������$�2d�A�000_°:��P(I$�����$��	@�,9NS��9NS��9NS��9NS��34'��W��BxȈ���`��P�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(*��#>*�)�r��A��62�2�	�Bj5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�� �z6c$ ��8r��)�#L鞎�� t���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� U�*�#�`p2@0Y�9NS��9NS��> `0� #8ļ�\�9/)��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4e�a��pX��9NS�����#�V��e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���̠3�H�GPy�r��)��`�3&d�2����������L�3Y��(
�#�TʙP �APg����9NS����c�9�3&dBA2d�����ɓ(�J&�Y��Id�A2d�����������������������������������������������������������������������������������������������������������������������������������������"B�$�I$_°:��P(I$�����*EH�a!�S��9NS�%�(<�9NS��9NS��9NSdd�М�^#	�"##��nf9@s�1s�1s�1s�1s�1s�13���������)�r��S����@����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N"�f2@ J|�)�r��A�3���>��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y���6"0 2!]p3ac<�L"f���:r��)�r��0���'ʜ����A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��`�d#8X�> g)�r��|�Fq
�	!�g�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�P�$2%\%�)�r����8G�A#����������	000
���6&~3� H�C
���	A���r��)�r��(,��<e��
�������2b��_
��|I$��	�&L�?�������������������������������������������������������������������������������������������������������������������������������������$�2d�A�I$����VAА
�$�@�?����Q(�O��4�3NS��9NQP����d��d�8Ld��i�9NS��9NS��9J��3�L3�x�1 ��2"129���9�c��9�c��9�c��9�c��9�c�� ��PU��F|T	�S��9J��)�`le e�@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'ѳ  %>Ô�9NS�,g�<���X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,lDc>��1
���y�r��)�|�f
�3A�8�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aі	�B)�`lr��)�r�2�*@hI�>��O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR ,�������9NS��QG����������@�$�H0�9R*EH� l!0L�`���9NS��9NS��9NP�|�xfLə$�@_����&L�Q(��f�I$000L�0�"x@�?�������������������������������������������������������������������������������������������������������������������������������������	L�2dɒI #Y���� R�"H$O���AА_��_ �3�S��9@`�d �$! �t*�<U�V�	���1���t�9NS��9NS��*�ϊ�0��W��BxȈ���`b�!�b�!�b�!�b�!�bg�AW71�P&9NS��*�����������@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j���D/C0T ���S��9A�i�3���>��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "��xaN3��9NS��b	�3 	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ,�S��ب> g)�r��̪����2� ��*�YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�P�$2%\%�)�r��Cc���001���������2f�Y���}>�O�����H��#��9NS��9NS��9NS��9NS4�3L��2��P+����dɊ±|+��D�Q2��dɄ	$O�������������������������������������������������������������������������������������������������������������������������������������D�	$I�e�f�X(
�#I$$O���5��f~3�APg�)�r��q2%\\r������Z��*؁�y��%�)�r��)�r��)�3�LgT$��nb"�D���nf9@s�1s�1s�13�������8f�)�r���3������`Nj5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�� �z6c$ ��8r��)��π�1��H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@ � f���S��9J����t@��B�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aњ)����P| �S��9M�U 4$�ɟEZ�=+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��y��� �����9NS�Ca}>�F?������$```R�#blM��C(�~? P
 A`�Y�r��)�r��)�r��)�r��)�r���:dc#
�@�P'����fY V��Y��I$���A �2aD���������������������������������������������������������������������������������������������������������������������������������������$�2fY�H�b�
�@�����"����/��Xe��f��i�r��(l�X#&|3� ,�e�, �WH�U�x�"��8�!P���`�dr��)�r��)�r��hN���W�nb2�Q��dnf9@s�1s�13�������8f�)�r��S����@����@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N"�f2@ J|�)�r���4Ό�$F@��X@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� 4��&pr��)�r��b�3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�4�pX��9NS�ٕQPB 3FA	,U��Q������O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI�� ��C"U�Py�r��)�!�0�>�O�������ɓ(�J!�!ʑR*F&& l&H�� ,��)�r��)�r��(<�3��d�RF@fRF@b�d�)�r��(J> �BL$�� H����L�1XV/�f�Y$�2��,�$	��������������������������������������������������������������������������������������������������������������������������������������D�	e�d����Y��
�@�P���@�?����/�a�2�Q�#�H�9NS�3���1��H,@Yb�X���nb�#�V�⬊� H���P���Py�r��)�r��)�r��g�@����UJ��,eY��@&F�c�1s�?�
���ϊ�1�r��)P| �8,�� ���j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�� �z6c$ ��8r��)��ρ��� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����fJ� �����g)�r��(��/0W#���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�3A�9~2g����)�r�2�*3���X�Z�=+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�Q��@g��ȕp�|�)�#L����8001����� H�dɚ�f�@�PG�?�����i��σ��9NS��9NS����t&/�)S��073�fg�@�(�̫�AL�S����9NS��> `l!&`j$O���&L��+°�_I #,�$fY  H�$O��������������������������������������������������������������������������������������������������������������������������������������2dɓ/��X
B�$�'������2�P�2D|��)�r��q�3�@�e�,@Yb�X����fJ���U�t*�<)�A�y� ���t�9NS��9NS��>�$g�@����U��Fi�xl 	��!�&
��A�a�r��)P| �8,�� ���j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�� �z6c$ ��8r��)��π�0���,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@$)S��S��9NQ�,^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4f�r�d��A�9NS��6eTT�ѐBK`�@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3�`� #1
�g�)�r��\������001����&L����(
6&�ؗ��$	BCc4�3NS��9NS��9NS����t��"4��B���&g��m5S����/2�e$d#L��r��(<� @a	0�P�"���2d�%��+ĒH�$	�&$H@�?�������������������������������������������������������������������������������������������������������������������������������������	$I2d̳,�000_°(
�#I$$O���/��Xe��d���9NS��	A��Xφy�� ,�e�,@Yb�X����p3`$)S?�$df�h�G�`�4Μ�)�r��)�r��A��1_�E*�Xq�2"�2"�gT$��2NS��9J��)�`le e�@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'ѳ  %>Ô�9NP�|�$FA U� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� � f��&i�r��)�3�e�����G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ����`N_����> g)�r���&2e��2� ��*�V���J�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI��@�g�P�$T�t*�(<�9NS���CO�с�����$ID�Q(
d̙�0�8�r�FA`�Y�r��)�r��)�r���d�`g��� W�\@���Du�{<�৒<��(!�@C����:r��)���x�P('����&L�Q(��f�I$e�	ɓ'�������������������������������������������������������������������������������������������������������������������������������������$H@�$ɓ$�@E�|+�@�B0$�@AD����D�}>�L�2G)�r��1�F�e���g�:@Yb�X���� ,�e�,@Yb��93�@�$)S1
�L"f��M���:r��)�r��)�r� �6bg
����l���r��)�r��g ���+� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���C4����ٌ� � ��r��(l�X# �*�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "�HR�#�	��)�r��8X��\�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h���ɟʃ�r��)�)�c&X�,2Ib�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI��@�g�P�$T�t*�0Y�9NS���CO�с�����&LB@I����8G��2�x��i�r��)�r��)�r��(<�3�1~	J��Ɂ�F��@�� м����H�S�
y#�D#@��A�� �,F�Ӕ�9J����x�P('����&LV��Y��I$���A �2�D�	�������������������������������������������������������������������������������������������������������������������������������������$ H�,�$I #Y��
�!��I	����$�#�p��$r��)��hXφy��fJ����� ,�e�,@Yb�X���� ,����3�71V@hȕr>g�8T#�3��9NS��9NS��9NS��9NS��*���/0W @Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'ѳ  %>Ô�9NPygFX# nb� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�����)�r��(��/0W&���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M*r2^R�d��A�9NS���1�,g��$�V
�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����U�j3�(���σ��9NQ!�1��}$�@_�$I$��F�؛�2�Q��~�C�`��|�)�r��)�r��(�'�� F|��B�a�fP����E0^��H�Q�)��S@��D#@��A�� �,�9NS�%� l"�@� H����L�2�D�+
��$�2��,�$	����������������������������������������������������������������������������������������������������������������������������������������&L�2��|+�@�B0(�J!D����I$G�2D|��)�r��qFFh&��� t���� ,�e�,@Yb�X���� ,�e�,@Yc#��g nb��%*b�#�U#�z3�c8���t�9NS��9NS��9NS��9NR����b�3rj5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�f�qp�1� S�9NS����t,�f*��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�@i�*���r��)�3�e�����G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��*r2^R�d��A�9NS�F��N2�xa�BK`���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�Z�=2��"�#�U	A���r��)�#�H�����%��ɓ$��A�!ʑR*F&& l&H�� X,T 3��9NS��9NS�F��N2O�)# 0H)��xS"�
+�O�<���L�H�S@��L���3(b0����9NS���@�P$O���$�Q(��f�I$e�	ɓ'�������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�I�f�P(!F�D H����I$���#�H��#��9NP,�����H,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@ 
����T�t*�|�Fp��y�r��)�r��)�r��)�r��g ���+��	�h0'5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�� �z6c$ ��8r��)��ρ��� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X� �� ȅtB 3M�US��9NQPU�f
�sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F���f2@�T��9NQN2�xa�BK`�@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI��@�g�e'�(�*b:P,��)�r��`����(

%���k
p�����3Fh�#�HF�Ӕ�9NS��9NS����tL�g�	�`�`��*��4/�C*b:�`��H�S�
!��04
`h��)��S@��S@�	���X<�3�)�r����@�P$O���&L�D�Q�b��Q(�&L H��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�H2���V�B��)J%�"���$�#�p��0Lr��)��#�q�g�<���X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���T�� t��Xe�"2��0Y�9NS��9NS��9NS��9Bp<�&�̌�L2 cP��@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��3A�8�8^��� )��)�r����e�"2�9e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����ИD�9NS��9E@yTHy��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F����* A�T��9NQN2�xa�BK`�@�g�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI��@�g�e'�`� #1
�l�S��9NQ!�1�2�Te��bbb~?�("��3�S��9NS��9NS����tA #>	3�0�0̠!��h��ʘB4
!����F�L�04
`h��)��S@��S@��eF pr��)��π<��@@�?����2e�DV��D�000e�d��"B���������������������������������������������������������������������������������������������������������������������������������������	L�3,�$�f�P(!F�D�2���```̙�2�1�r��(l��d��g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���G3�L�g�:X�,2��#�	� �f��9NS��9NS��9NP��8,��9�	!p��h0'5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�h0'ѳ  %>Ô�9NPygFX# �*�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb���*�A �#�z3�S��9NQ�,^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���iS���1� ����)�r�p�ɖ3���X�Z�=+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'���A����T6G)�r��)�*
�8��r2d�����t�9NS��9NS��9NPM3��# 8?�_����"�W��#��؄h�G��F�D#@��L�04
`h��)��S@��L���3(b�=2`�4Μ�)�r��x(
	�'�����(�J"�|_J%���dɄ	���������������������������������������������������������������������������������������������������������������������������������������2dɓ/��X
B�D�Q&L����&L��3&d��r2r��)�� 8�"�K�6�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
��K�e�2��|A3�,��)�r��)�r��)�T�J��&��$|�X&1�f�p cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@ơ�	�A��3@	O�p�9NS�F�і�� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X������>g�8�9NS���P^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���iS����P
��r��)�2A4L�x6"1V���J�O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����lD`��d�h<�9NS��9NS��9NS��9NS��9A�i�	��JT�L��ي��xB�j2�04
y#�O$x)��Q�(�hB4
`h��)��S@��L�04
`h��)��Q�)��PC2��# 89NS��*� ��P('����&L�Q(��f��D�e�	ɓ&L�'�������������������������������������������������������������������������������������������������������������������������������������	$H@�$�A�I$����V�B��|_
�D����A �*EH��0Lr��)�� 8�":h@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �WL�g�:X�,��1���t�9NS��9NS��9O��� �Pٌ� �O�Hx��!����j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1�D/F�d� ��S��9@`�d2��W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��`�� � f���S��9NQPU�f
�sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�9/)�  �*��r��(��x2��� ��e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�@g���Dd6G)�r��)�r��)�r��)�r���4΄��%*��*�@�=P�H�)��`h�G��H�S@��L�04
`h��)��S@��L�04
`h��)��S@��S@��ee$dr��)��π<�L$�� H����$ID�Q�b��Q(�fY  H�$O������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�I��
�!��/�`�"��� �e��2fJ�W#')�r���4΁�<��^A��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��`�� 2!]3�@�c<�̐��y�r��)�r��)�r���P_��^͘�  p��x��`�d @Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�A��l�H 	O�p�9NS�F�і�� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���G3�A 4��&pr��)�r���2�2�qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��*r2^Q�* A�T��9NQ�	��VE[&�@F+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'���A��U�y��r��)�r��)�r��)�r���4Ίq�|I��/�~^Ȭ���Du�{��F�D#@��S@��L�04
`h��)��S@��L�04
`h��)��S@��D#@��A�� �,F�Ӕ�9NP6@�P$O���$�Q(�±|Q(�L�A �2aD��������������������������������������������������������������������������������������������������������������������������������������@�!D�	Y$�/��XB@�!��$O���&L�R*EHCar��)�� 8�"�K�6�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���G3�@��XX�,���4Μ�)�r��)�r��)�r�A~���  ��2�2� cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j5�A��l�H 	O�p�9NS�%�,	�@q�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��̕@ � f��=�)�r��(�*��3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�J����f
�`�*��r��(��x�"��`� #����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�`� #�� t����<� �qr��)�r��)�r��)�#L�L_�R�=2`ng&�U�S���&}�iE0^�$x)�<���Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��D#@��PC2��# 8��t�9NS� M�P(	�����(�J&�Y��Q(�&L H���������������������������������������������������������������������������������������������������������������������������������������D�	Y$�/��XB@�!��L�?���L�2�T�� ��9NS�F��8�":h@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����We�"2�#��9NS��9NS��9NS��	O�p'��  ����/0W @ơ�	�h0'5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j���D/F�d� ��S��9A�i�`H�� ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� 4����9NS��9E@yT��+��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=T�d��0T�P_�S��9FH&��Yl@����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�Z�=*�5�YI�d��X/32U䗐l"��� OM�`�	��J>S��9NS��9NS���$�2�2*�!�f�1�g�D���/f�O$x)�04
`h��(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�)��PC2��# 8��t�9NR����xa&�D�����"J%��_��D```�2aD�	�������������������������������������������������������������������������������������������������������������������������������������$�2d�A�000_°(
�#����'���ɓ&*�P� �0�9NS�%�df�i
� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�d�h<�9NS��9NS��9NS��9NS��*���1����'̤ ��e�a���`Nj5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��"�f2@ J|�)�r��(<�`H�� ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� 	J�&3NS��9NQ�,^`�M�M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4���y@�1>
��r��)�2A4*ȫb� ��e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?����TЫ@�#�U	�L�P���S��9NS��9NS��9E8�>������? �,���'���)��y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
`h̠!���S��9BPy� �&�a&�D����dɔJ%XV/�%��H$&L H�$O�������������������������������������������������������������������������������������������������������������������������������������D�&L�2d�H�/�`t	�`_±2d����2d��x�`J>S��9Ba4��Z�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e���X� ��M��)�r��)P| ʃ�r��)�r��)�r��%>��3�b3@0 �32e e�,��j5���@@Ơ cP1��j5���@@Ơ cP1��j5���@@Ơ cP�8^�`�)��)�r��f�e�"2�9e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�y����%*b> ���r��)�3�e�� ��sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F���3�O����)�r��M��*؁6"1YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR$�V����f*��x`�1L�6G)�r��)�r��)�r��(L_�PH)�D^e\�6������F�O$x)���04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
`h̠!����i�9NS�� @a
D����dɔJ%XV/�%����2d����������������������������������������������������������������������������������������������������������������������������������������	$I2d̳,�000+
��:��B05��dɓ����ɓB�U `T 3��9BPy���t*�<��`��e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�S��L�9NS��6FL��Q�e!A���T 3��9NS��9NS��> a)��x��M���1�f�p cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��j��  %>Ô�9NPygFX# �*�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb���*�HR�#�	��)�r��8X��\�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�Рp Fq��T��9NQ�	���� ��e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'�BK`�<��/ �EYl@��<�
p�ɀ�f��9NS��9NS��9NS��9E8�>��E�&�C*a�)�<�৒<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L���F�A�� �,F�Ӕ�9J�� �&�a&�D�����"J%��_��D```�2�D��������������������������������������������������������������������������������������������������������������������������������������@�!D�fY ```�Q(��f�B0/��X�2����2dvG`���xJ>S��9Ba4 ���,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���nb�
EB>9NS��9Bq��M����Wpl4�dA���T 3��9NS��9NS��	O�p'��� ��l�ɔ����L2 cP1��j5���@@Ơ cP1��j5���@@Ơ cP1��"�f2@ J|�)�r���4Ό�$FA U� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����/32U ��G�89NS��9Fp�x���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѡ@�( ���/�)�r��0Y�
M���VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�Z�=+)?���͂�� �WA 	J�dJ�L"f�p�Ƀ��:r��)�r��)�r��)�r��)�T�L̠!��)��y#�O$x(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h̠!����i�9NS�%� l!&`j$O���&L�D�Q5��e�D�$	�&$H@�!D�������������������������������������������������������������������������������������������������������������������������������������$H@�$ɓ$��D�k5��@�Q|_
�ɓ����D�bl@�<	A���r���4΄�&i
�29�&r@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���G3�B��P���S��9J��f���{3$���1*@��x# ns4�dA���T 3��9NS��9NS��	O�pT�@�"	�3" �z5���@@Ơ cP1��j5���@@Ơ cP1��j5�`N"�f2@ J|�)�r��(<�`H�� ��@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd� 4��&pr��)�r��b�3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�B��P�'�P_�S��9@`�d� ����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�h��$�ɟF�@F3�@�c<�X�����͑�r��)�r��)�r��)�r��)�r���:	3���"`h�G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
y#�D#@�	��S��0ygNS��9@�<
D�����"J%��+��D```�2aD��������������������������������������������������������������������������������������������������������������������������������������$�2d�A�I$��f�X:������'�����6&�؁�xT 3��9BPy�G��gЫ@�#��g$� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �WB���	���9NR�����"T�R/F��( T2� N^ Џ�79�n2 �pA>�$�9NS��9NS��*�J|��<� �13�$+�8^�X&1��j5���@@Ơ cP1��j5���C4����ٌ� � ��r��(J>X# �*�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yc(�/32U ����)�r��(��/0W#���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4(
s`��8r��)�2A4� ����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR6"1e��/ �@�/ p2B�&2a(<�9NS��9NS��9NS��*��T����)�r��(�'��r�+�O�F�O$x)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��<B4
G� �G	�)�r��A���<P(	�����(�J"��_J%,�H&L�@�!D��������������������������������������������������������������������������������������������������������������������������������������@�$ɓ$�@E�|+��H/��X�2��� H�blM����4Μ�)�r��=���ds0L䀲�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��	�p3��4Μ�)�T 34�dJ��E���y�e!���nx<�"�d�AxB<F@��8�����p�> g)�r��)�r��)P| �S��P)̀g�HW�p��L2 cP1��j5���@@Ơ cP1��j���D/F�d� ��S��9BPy�2��W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��`�� � f���S��9J��3�e���ɸ�)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F���aNl ��S��9@`�d� ����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?�����O�e'���!%��lDb�3%PGB�ʘ��T���� ���t�9NS��9NS��9J��|�ɑ��S��ؿ3�N���/�)�r��(<�3�ng&�W��<�৒<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��R< zT�LF�Ӕ�9BPy� �&�(
�����D�J%Y��Q(�F	�&$O���������������������������������������������������������������������������������������������������������������������������������������"I�&H$d�H�/�`t	�|+&O����	lM�� @a	A���r��)3ќ	 JT�G3�H,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r� �f���SH��&�ɹ��nx<��2����y EP�N "���x����q��#A4*�P| �S��9NS��9J��F�\g � �bg�HW�p��L2 cP1��j�����@@Ơ cP1�f�qp��PS�9NS����te�"2�9e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,����3�A �#�	��)�r��8X��\�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�Рp)̀� ��r��(��xS��lDb���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����VR+)?���͂��g�<���x`�1�*��g��4Μ�)�r��)�r��)P| �S�	��:3@0g�HWі	�B3A�9��!_E@yT��9NS�6@ng&�W��<�৒<��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S�
!#� g����ygNS��9@�<
D�����"J%��+��D�$�,�$O���������������������������������������������������������������������������������������������������������������������������������������"B�&L����D�Q5��b��_&O����	d�z @a	A���r��A�#�	�@�1e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��U�O��G�g)�r��A�3M�D���^���s����y7<M��s�����t�d6B/)S����	�zeg1V����9NS��9NS��*�|qN`aNl=2B�����f�
f3A�8��4����@@Ơ cP1��"�f2@ J|�)�r���4Ό�$FA U� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���P�$^fd� 	J�&3NS��9NQ�,^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���hP8
��	O�p�9NS�6ELGB�lDb���YI����VR+)?�����O�e'��YI����VR+)?�����O�e'��YI����2Ib�X��Z��*؁=7��&2`0Y�9NS��9NS��9NS��> c>l�N`aNl�3r3A�8UJ�9���F����*��/�)�r���d� ng&�W����H�S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x(�h���9���t�9NR����x(
�����ɓ(�J"��_J%���dɄ	��������������������������������������������������������������������������������������������������������������������������������������D�dɓ&L```�Q(��f�I$L�?���́�/E�	A���r��)�*�� � f��9 ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y`71V?�"���)�r�����7�f0I��&�ɹ��nx<��&�ɹ��nx<�� t�d EP�N "���x ���T�XF�h8T 3��9NS��9NS��> c>l�N`aNl=2B�����f�
f3A�81��j5���B �z6c$ ��8r��)�#L��Dd��U�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����fJ�B 3H��g)�r��(��/0W#���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�J���9�S�9NS��	A���Dd� ��e'��YI����VR+)?�����O�e'��YI����VR+)?���ʴFzVR6"0��d`HR�*b:P8�!P����i�9NS��9NS��9NS�%>�&F��f2@ /�>e e�@�(�A��F�z4sѣ��6�_�aNl ��S��9A�i�?�_�+��)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��(�h���"��i�9NS�%� x���"���2d�%��+��D```�2�D�	��������������������������������������������������������������������������������������������������������������������������������������D�	L�1����D�_±$�&L�����&`jX�`�|�)�r�p�ɂ@i���3��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����p3`S��*��r��)P| ��q�*b��s����y7<M��s����y7<M��s����y7<M��U�^��	3=	!T�O	�R��p�> g)�r��)�r��)P| �|�"���zd�}�1��j5���B �z6c$ ��8r��)�#L��Dd\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�3%P! �|A3���9NS�g ���+�qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��
@�)��)�r����e�"2lDb���YI����VR+)?�����O�e'��YI����U�j3ҭQ������O��@Fp3ac<�XٕQP6G)�r��)�r��)�r��%>���0T	�3#,�*�S�h�G=9���F�z4sѠ	U*�0�6 ϛ!�9NS�F�����B���H�S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x(�h���"�S��9NP<��A2d����@�%�DV/��D�000L�0�"���������������������������������������������������������������������������������������������������������������������������������������"I�&000I$����V(�J$ɓ������X�`ygNS����tS��LB 3L�f	��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]
E8Ld�S��9J��f���SH��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��*�@*q�4#�'�ʨ��3�fT 3��9NS��9NS��> di�U�8,��9�	 �"� cQS������B �z����8r��)��!��� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X�<��̕@ � f��&i�r��)�3�e�����G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��
@�)��)�r����e�"2lDb���YI����VR+)?�����O�e'��YI����VR$�V,^Iy�*ȫb�HS��L%�)�r��)�r��)�r�A~�d ��`aNl�3rT�d��	U*��G=9���F�z4sѣ���h�@�U0aNl�6B	�r��(<�3����"�p"y#�O$x)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��<B4
G� �G	��4Μ�)�T 06@�P$O���&L�D�Q5��e�D�$	�&L�>$O������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000I$��f�YD�Q2̲G���$$�LK,|�I�r��(�	�� � f��9 ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�� ��|r��)�T 34�dK٘�&nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��l �^R�f0I�R��q��6FL�9NS��9NS��9NS�/�>l�Nb�f�K��Ȉ8^���C4�Hy~2g��/�)�r���4Ό�$FA U� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����/32U ��L��)�r��(��/0W&���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G= �R��
s`��W9NS��	A���Dd� ��e'��YI����VR+)?�����O�e'���A���X	 JT�C"U�a4T#�0ygNS��9NS��9NS��>
��	@3f2@ /�>"��pn �h�G=9���F�z4sѣ���h�G=9��a*����#O��r��)�#L��r��\�H�S�
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)���� 3��Bp<�3�)�r������	05'����	Q(�EaX�(�J#Y�H'�	��������������������������������������������������������������������������������������������������������������������������������������ɓ&L� �e�I "���%�2d����
�����)�#L�	�� � f��9 ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y`71V?�"���)�r� �f���{3$���:P2�&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��R�LU"�g�$*��?  YU6FL�9NS��9NS��9NS�/�0�/�L�U��h�#��e e�p��N�Ҡ���)�r���:2��W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�@g��y�����> ���r��)P| �p�x���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѠ	U*�/�>3��A9NS��	A���Dd� ��e'��YI����VR+)?����H|��lDc>��3�� e����g$A�)�r��)�r��)�r��%>�PU g���f�
f�=9���F�z4sѣ���h�G=9���F�z4sѣ�� J�T��~	�6B	�r��(<�3����"�p"`h�G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
y#�O$x)=D'��:r��)� �&�(
�����D�J%XV/�%��H$&L H���������������������������������������������������������������������������������������������������������������������������������������D�	L�1���I$_±D�Q&L������@�~?�`���9NQN2�xb�3%P@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���nb�
EB>9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��l �^R�*�zM��0� q��6Fpl�S��9NS��9NS��*�% �8,��� 8X�*��r��)�#L��Dd��U�� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����fJ�B 3H��g)�r��(�*��3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U08_�|g͐�r��)��ρ���e��O�e'��YI����2Ib���*��K�6VE['��0S��LF�Ӕ�9NS��9NS��9J��3��A�2������	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�p��ϛ!�9NS�F�����B�04
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�F�O$x(�h���9���t�9NS� M�P(	�����(�J&�Y��Q(�&L H��������������������������������������������������������������������������������������������������������������������������������������� H�dɒ	Y$�/��X�Q(�fY#����@�~?�`�Y�r��(�	��c<�y���2��"�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���nb�
EB>9NS��>�$�7�*�z7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��a"�1T�Ђl�6e��*�&�ə�)�r��)�r��)�T 3�/�A�9NS��9NPygFX# nb� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X����/32U ��G�89NS��*��*��3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U2�f�F|�')�r��)�� D+�$>L�+)?���͂��^fd��U�xS��������:r��)�r��)�r��)�T�&F���d��p���8^���Q��)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�p��ϛ!�9NS�F�����B�04
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�F�D#@��R< z8�N9NS��*���&`j$O���$�Q(���|Q(�F	�&$H@�?���������������������������������������������������������������������������������������������������������������������������������������&L����$�b��Q(�&O����@�~?�`�Y�r��(�G�e��2�nb� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�� ��|r��)�T 34�dJ��E���y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���A��4�"	�B|ٖ/�,���#86g)�r��)�r��)�r��)�r��(J>X# nb� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���P�$@Y`A �#�z3�Py�r��)�3�e�� ��sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�FL�\��NS��9NSfUEB�28ds0L��<���XX�,�6eTT�͐<�3�)�r��)�r��)�T 0��p<��P��f�sa*��7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U08_�|g͐�r��)�#L��r��\�F�O$x)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��<�G��� 3��Bp<�3�)�r���� M�$�LB�����ɓ(�J"��_J%,�H&L�@�< H��������������������������������������������������������������������������������������������������������������������������������������$�2d�A�I �aX�/��X�2����
�����S��9EB>,g��p3ae�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "Ч�S��L�9NS��> fi�ȕ1T�ѹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ�� ���ĩq�G��!>l��UDO�x�9NS��9NS��9NS��9NS�%� ``71VX���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�XB 3H�����|�)�r��b�3r9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U22f��g͐�r��)�r����ٕQPe�"22%\�HS��L6G)�r��)�r��)�r��g͐�3�e��9����S���%T�c���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�S��'�|�')�r���4Ο�/�����h�G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��� 3ҧ=2`�4Μ�)�r��x(
�����ɓ(�J"��_J%���dɄ	�������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000I ���V/��X�H2����1?��`�Y�r��(�G�`tʗ� dB�lDb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���nb�
EB>9NS��*��n2%��`�7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q� �	�B|ٖ/�,��� �r��)�r��)�r��)�r���:�W���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��@i3ќr��)�r��b�3rn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѠ	U*�W3M�>l���9NS����t6@0Y���t�9NS��9NS��9NS�/�L�/f�d� 8_�|�@�ʜ����A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��O���NS��9A�i�����m04
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�<���R< z8�N	A���r��A� @a
D�����"J%��_��D```�2�D���������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$�|_
°�_	_����!̩�2��X,�9NS�T#�0:eK����,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r�����7�f0I�"�ds����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s��J�'# A�
�˃`2���Q�2NS��9NS��9NS����t&3J��� 
��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�@g��e� 4����9NS��9Fp�x���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѡ@�( ����S��9NS��9NS��9NS��9NS��> a)��x��M��`�d 	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��O��P�9NS���������S�
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)���� 3��Bq�r��(J> �BL$�� H����L�2�D�k5��%��H$&L H��"B����������������������������������������������������������������������������������������������������������������������������������������"L�,�000I ���V/��X�H2����1eL����g)�r�����*^ ��X@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt)�A �9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d7<Hĩr0�Fi�ȃ�������9NS��9NS���͐L"f�?� ��L�9y��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y` dB�	 JT�|�Fq�r��)�*ʠ��\�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�8^�p�P| �S��9NS��9NS��9NS��9O�����Fp�0�6 �#��T�d�����z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G= �R�����>l���9NPygA �p)�X04
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
!#� g�����9NS���@�P$O���$�
±|Q(�F	�&$O��������������������������������������������������������������������������������������������������������������������������������������$I2d�	  |_
��|+	_����!̩�2��X,�9NS�d�h<�R��f*�(� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �WB��N3��9NR�����"^��	3s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y#�	��g�8@e��"F�h8|�I�r��)�r��)�#L���xL"f�?� ��L�f*��3%P@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb� "�A �#�z3�S��9NQPU�f
�sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�� ����S��9NS��9NS��9NS��>
��	@2�d��p���8^������A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qS@�~	�J��)�r���S8Ȭ�<���L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�Q�)=D'��:r��)P| ��<
D�����"J%���k(�J&Y �L�0�"B���������������������������������������������������������������������������������������������������������������������������������������	$H@�$ɓ$�@B��_�f�A �����0�9�2�T�3LӔ�9NQ�	��:eK����,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��U�O���y�r��)�&i�ȗ�1�L��y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��U�F%H�� �d����)�')�r��)�r��)�#L�G�a0��� �Ы@�71V�9 ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+���LG��g�)�r���<�� ��sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)�NFK�e e�g���J��r��)�r��)�r��)P| ʃ�� �N�ј*�=2B���aL̈́����A��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�SM�����r��)�	3���@��Q�)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S�
!#� g�����9NP�|  	����"���@�%�DV��D�000L�0�"���������������������������������������������������������������������������������������������������������������������������������������"I�&000I �aX��b��H2����� �3��*��9NQ�	��:eK����,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�"���)�r� �f���SH��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� � ��P �'�q��>�$�9NS��9NS��9NPygEB>##4B��:h�f*��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Y`HR�#�z3�Py�r��)�*ʠ��\�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�S���@��	 g��`��
��r��)�r��)�r��)P| �|�"�������	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�SM��2di{9NS����t
g��S@��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�H�R< z8�N��t�9NS���@�P$O���$�Q(��f�He�	Y�H'��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�H2�$�|_
ƳY��H2�����# 0�*
�8�9NS�d�h<�R��f*��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� D+�O��G�g)�r��A�3M�D���^���s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q�78<NS��9NS��9NS��9NS�T#�08�!VE[$t*�<��U��fJ����� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��f	��@iL��9NS���2��f
�sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSB��P�8^�ffF`�8BS�*��r��)�r��)�r���*�#Kٳ  ��2�2�p9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�l�ɓ#K��r��(<�3��S8Ȭ���04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
y#�D#@�x@���L�<�3�)�r����@�P$O���&L�D�Q�b��Q(�&L H��"������������������������������������������������������������������������������������������������������������������������������������� H��"I�&000I$����V�b�``c����P( ��APg�)�r��f�U�V�����3�H���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]
EB>9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d EP�`3��*b�*��r��)�r��)�r��)�r���:*���dU�GB����X@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��`�� � f���S��9NQ�,^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�n �iS���Hx/�>_����g�P_�S��9NS��9NS��9J��2F|�F`�	�3#4S3a*��7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���&�̙24���)�r���S8<�x04
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��F�H����!8F�Ӕ�9BPy���x�P('����&L�Q(��f��D�000L�0�"x@�?�������������������������������������������������������������������������������������������������������������������������������������$I2d�
%�|_
ƳY�``c����P( ��APg�)�r��f�)�AW���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��*��r��)P| ��q�/fc����nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��{3$͙b�#&f��)�r��)P| �S��9NS��9NP�|
�|FFh&��*؁/$��ap3a���3��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�3%P! �|�Fq�r��)�3�e�����G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G= �R���`N H��aNl�,3��A*�P| �S��9NS��9NS��9NS&F��8_�|���y@�U1�F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4A6fdɑ���9NS������E`��(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��(�h���"�S��9NP<��A2d����@�$��k5�J%���dɄ	�������������������������������������������������������������������������������������������������������������������������������������� H��"I�&H$d�H�k5��f�����"���:��4�3NS��9@`�d� �������� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��)�c&r��)��σ4�dK٘�& �����s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q2��6FL�9NS��9Af�@�͘�6FL�*��r��)�r��)P| �Py�)�c& �$*ȫb�������TX���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�3%P! �|�Fq�r��)�3�e���ɸ�)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��X&�l�ɳ  d�����8T 3��9NS��9NS��9NS��9J��3�e�A��n �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�ٙ�&F����9NPygL�*
dVL�F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��O$x(�h���"��i�9NS��> `l"�@� H����L�2�D�k5��  ���2d��'��������������������������������������������������������������������������������������������������������������������������������������@�$ɓ$�I$k5��f�X��������:�����3LӔ�9NP,��$FL�g�:@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt)�A �9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ ����r��)�%��W��2"�+�b8W�dd�Ӕ�9NS��9NS��	A���	����*�#�e䗐l  ȅt���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��3�H���T@�1L��9NS���P^`�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ�����) #/��'��?�24��A~*��r��)�r��)�r��)�r��)�T 1Na�	�Bn �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4*�SM��2di{9NS����tq�)�X04
y#�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�<���R< z8�N��t�9NP�|�xa&�D����dɔJ%Y��I ��A �2aD��������������������������������������������������������������������������������������������������������������������������������������$ H�dɒ	YD�Q/��X�k5�	�����t$��f��)�r���4΄�&ic<�y��� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�, �WB���	���9NR�����"T�R/F�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%��`��� l���r��)�|�H�#���|���|���q^#¼ ��8f�)�r��)�r��(l��U�pp�R�^Iy� �WH,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb���*�HR�	�LӔ�9NS�T�Ax���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G= �R���aL���
� Fq����ϛ!�> g)�r��)�r��)�r����	�`���$�#��9NS��> c8XD/F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�MM��2di{*��r���4Ύ"�\@��S��G��04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��� 3��Bp<�3�)�r��l"�@� H����$I$5��d�```�2aD���������������������������������������������������������������������������������������������������������������������������������������D�&L```�Q(���k5��?���AА_��_�i�f��)�r��$A��0��X\r�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X ��?�#$A�)�r���<d���"^��	3s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���f0I��� 6Fpl�S��9O�x��`_�129���nf9@/3�D'��W��p8^�М3S��9NS��9NS�%�̪��`b�28^Iy� �WK�̕Ae�,@Yb�X���� ,�e�,@Yb�X���� ,� 2!]��> ���r��)�*ʠ�@��=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M
C4S1ٙ��* @N���/�A�9NS��9NS��9NPygL�2@x�S*eK���������X,r��)�T 1PU �z�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�ٙ�&F����9NS�q��"���)�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��F�H���S��0ygNS��9@�E�@@�?����2d��k5�@@!���dɄ	����������������������������������������������������������������������������������������������������������������������������������������	L�2dɒ	Y$�5��`�:�����Y���~6�#�H�9NS��9@`�d����� H�U�x���,@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e��
�S��*��r��)�&i�ȕ1T�ѹ��@�Cs����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q�� 6FL�9NS��>�$/fT�@ !�C�1�C73����"�D�*6b�34�9NS��9NS��9@`�dlʨ��*�#�f|3�29�&r@Yb�X���� ,�e�,@Yb�X���� ,�e�,! �|A3���9NS�T�Ax���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�Aҧ#%��/�>_����g�P_���r��)�r��)�r���X,��r28㘘��"�T�!HR(�J �P(e��!�0�9NS����tg ����sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSDffFHϑ��r��)�8�NXqGQL��
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)���� 3��Bq�r��)P| ��<	0�P�"���2d�  ��k$��Cɓ$ H��������������������������������������������������������������������������������������������������������������������������������������$ H�dɌI #Y���� �I���+��#�p&	�c��9NS��9A�i���H��X���� ��X���� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd���P���S��9J��f���SH��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��1�Lf��3�fr��)�|�H�#������1�C�1�C�3s1� yy�%�dE\f��f�@�#&f��)�r��)�r��(l��U 2��Xdpφy��fJ����� ,�e�,@Yb�X���� ,�e�, �WA 4&3NS��9NQ�,e e㞍�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G= �R���`N H�! �b3�e�|�%A�9NS��9NS��9NP�|
����C@�$2�P�6&�؂�@�����"y2d�P�@l')�r��(��Ѹ�)����z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���i��)���I�1]9NS��9L�*,��#������F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�(�h���"��i�9NS�F��6@�P$O���&L�D�Q5��d�```�2aD���������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$���kAАI$�������Y �lM��q�`�Y�r��)�r��(l��U 2�Ō�2�|3�29�&r@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�X��� ȅt)�A�F�Ӕ�9BPy�f���{3$���s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<K٘�&3� �34�9NS�����F�##��9�c��9�c��9�b�2	��!���L�	��xWٕ	��{>�$�9NS��9NS��9@`�dlʨ��,g��3�@�y��� ,�e�,@Yb�X���� ,�e�,^fd� 4����9NS��9Fp�x���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�B��P��!M��6c$ �x	O�p�> g)�r��)�r��)�T 34�3@�< @��3&dP(�f�d���2d͉�6%�*��r��(���8^��M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"� H�����4Μ�)�r�TXq`h�G��F�D#@��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��(�h�G��� 3��Bp<�3�)�r��l!&`j$O���&L�D�Q5��d�```�2aD�	��������������������������������������������������������������������������������������������������������������������������������������D�	L�2A �$�@F�Y�BAD�Q'����Y��G�,X��#�H�9NS��9NS�� �	�LҦ#�U#�V��nb� ,�e�,@Yb�X���� ,�e�,@Yb�X���� ,�e�,^fd���P���S��9J��f���SH��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��1�L ��dg��9NS��34W���2�1�C�1�C�1�C�1�C�0���2;L�U��F�	��{>�$�9NS��9NS��9@c8�#�z3��D��3���� t���TX���� ,�e�,@Yb�X ��@i3ќr��)�r��b�3rn �h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���9/)��������ɟ̙^ς����9NS��9NS��9@`�d�1bŌLLJ�R*E�@�Q(�	���&L��X�c��9NS�g �tD/F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M/0W!8NS��9NS#
��. H�)��!��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�(�h���9�	A���r��( �I���	���ɓ&I �f�YD�Q&L�@�< H��������������������������������������������������������������������������������������������������������������������������������������$�2d�A�I$��f�X(
/��X�2����	k5��P�D �0Tq�r��)�r��)�*�̐�"���K�6 dB�@Yb�X���� ,�e�,@Yb�X���� ,�e�,@Yb�3%PL�x�1�9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ �ə�)�r���ə��F  ��P9�c��9�c��9�c��9�c��9�c��9�f�`�dv �ȫC0��6b�����9NS��9NS����4����`H��3���� t��`��e��3�H���� ,�e�,^fd� 4&3NS��9NQ�,^`�G=9���F�z4sѣ���h�G=9���F�z4�A�a*�����@��B���2�>l�����)�r��)�r��)�*
�8�Q~?�P�F�؛P(e�	����2f@��ŋ�)�r��8XD/F���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M$|HN�Ӕ�9NS���B�"���@��Q�(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L���F�H���S��0ygNS��*� �I���	���ɓ&I �f�Y$&L�@�?��������������������������������������������������������������������������������������������������������������������������������������@�$ɓ$�I$k5��@�Q��k$�����@�$ɓ1fLə?���C`X,r��)�r��)�#L�	��X��Xφy��fJ����� ,�e�,@Yb�X���� ,�e�,@Yb� "�VE[&̪��)�r��A�3M�D���f�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%��`� !<@���9NS��6FL��1 �a �L�1s�1s�1s�1s�1s�1s�1�`��L���Ȋ��/ l6b�����9NS��9NS���͑3ќT�t*���Lg�<���3%P@Yb�X����/32U ��lʨ�r��)�r��b�3r9���F�z4sѣ���h�G=9���F��"��X&	��!_F`��^ς����9NS��9NS��9A`�Y�#�H��*eL�#�pP(J%dɄ	����2d́�/@�$	�)�r��8+�R F^n �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�G�$��x��t�9NS�q��"����/b�Q�(�hB4
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L���3(b�=2`�4Μ�)�#L���@��d������"J%���k(�J#ɓ'��������������������������������������������������������������������������������������������������������������������������������������$�2d�A�I$����VAА�� �Q(�	�����D�I !@�P}>�K,d���	A���r��)�r��(l�����!�*�t*�<��U�G3�H,@Yb�X���� ,�e�,@Yb�X����fJ��R�)�c&r��)�|�I�n2%��`�7<@�@�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%��`��� l���r��)�l���+�b� �b�!�b�!�b�!�b�!�b�!�b�!�b�!�bg�A{ ��&r*ђ/ l6b�����9NS��9NS�F���#Ba4���UA 	J�\s#��g$� ,�e��̕@ � f��&i�r��)�*ʠ��\�z4sѣ���h�G=9���F��"��� ����/�L�	@3�/�A�9NS��9NS��9NPX,d���q�LLA�x)
B�D�Q&L������də ^�,#L��r��(��1/0W&���z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�M�M$|HN�Ӕ�9NS���L�=04
!��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
!������ �� g�S��9NP ͉�6$ɓ����D�J%XV/�  ���2d��'��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�I���� B�f�Y2d�������L�3Y��lM��111��<Tq�r��)�r��(<�3�$A�p2AO�	
�p3ae�,@Yb�X���� ,�e�,@Yb���*�:eK��	���r��)P| ��q�*b��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���f0I��� 6Fpl�S��9M��3Ex�@ �@ !�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(���U*�3�"���f O�x�9NS��9NS��9A�i� �	�L�!�*���L�9���3�� "Ҭ28lʨ�r��)�r���$|��M�h�G=9���F�%T�c4���S� g ���W*��r��)�r��)�r���X,�Q~?����6&�
	������də ^� H9NS��9FHϑ�x��7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�#�Bp<��)�r��Nzd�3�:�`��F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��Q�(�h��(�E`�9~�͑�r��)��`�6&ę2����2d�V��D�000L�0�"x@�?�������������������������������������������������������������������������������������������������������������������������������������$I2dɓ&000Q(�A�t$
B��)
B�D�Q'������ɓ�!H�"�eL�� �0��)�r��)�r���:)�c&zn3�e��g�:@Yb�X���� ,�e�,@Yb�X ���*^8Ld�S��9O�x�3M�D���^���s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<K٘�&3� �34�9NS��34W���2�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�⁚_�R�9~=�l�	P| �S��9NS��9NPygFH&��a4���UA 4����B 3L�pp3�Ӕ�9NS��`p��UJ�9���F�z4�J��A�� �323@0��t%> ���)�r��)�r��)�d�����<ʙS*dC.��(
f�Y2d�������$$�LO����r��)�2F|�K��ɸ�)����h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�>$'���r��)�T�L@A3=04
!04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��S@��S�
!04
+�O�� 3�73�f���9NS��9@06&�ؓ&O����	Q(�Mf�YD�Q&L�@�?��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�Q(��f�B0�!H
	_������"��@�}>����U��P| �S��9NS��9@`�dlʨ�2%\B 3L�g�:ds0L䀲�� ,�e�,@Yb�X���T
�*؁�1�9NS��*��n2%��`�7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y*q�� 6Fpl�S��9M��3Ex�@ �@ !�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C L�(���U*�3���_�f�@���9NS��9NS��9FH&��a4��f��	�$A�)�r��)�|�S���@��B���f�s) #/��'��?�24��A~9NS��9NS��9NS��r�FK,bbbT��R1Q(�B����������"E�A��~9NS��9FHϑ�x��7E4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=n �h�#��3�b�r��)�r�9�L�H�)��!��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��)��Q�(�h�G��F�H�)���\�� 3�? �@�	��Jr��)�r��(��F�؛d�����dɔJ%Y��I �	�&L�?�������������������������������������������������������������������������������������������������������������������������������������� H��"I�&H$d�H�k5��@��␤)J%�"����ɓ(�J%�|+&O��"I  �2迋����L�2A(<�9NS��9NS���$�	�LЧ���Z������`��e�,@Yb�X���G3�EYl@�p�ɜ�)�r���7�*�z7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y/fc��? dd�Ӕ�9NSdd��^# L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�0�⁖2�,�����U	()���x�9NS��9NS��9A�i���t�9NS��9NS��>
��3�e�`� �1�2�i�Uʃ�r��)�r��)�r��(<�3L�4Ca~?�P�F�؛t	Y �$O��������L�2�@�~?�S��9NQ�3�b^`�M�M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�^`�Fp��r��)�T�L@A3=04
!��F�D#@��L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h�G��H�S�
`h���/`�m3(`0�0q���F�Ӕ�9NS��9NP<́�/Dɓ����ɓ(�J&�Y��&L H��"B���������������������������������������������������������������������������������������������������������������������������������������$I2d��,�I��
�C�B��_°@�?����H(
��6%�G�ɓ&�� ��� �3��`�X,�9NS��9NS�F��P����d��e��/ �@�
�e�,@Yb�X��`�ȫ"��N3��9NR�����"^��	3s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���@�? dg��9NS��34W�� ?�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���&�2���U*�3���_�|T	�S��9NS��9NS��9NS��9NS��9J��|��*�P| ʃ�r��)�r��)�r�����3L�<̩�2�D2�ˢ�@��k5�&O����������	(
����r��)�2F|�D	 �n �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦR F^3�e�S��9NR�=2`�. L�F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`h��(�hB4
y#�L�5S&�(�̫��/�`b�d� �4Μ�)�r��)�r��i�f����������&L��f�I$H$dɓ'��������������������������������������������������������������������������������������������������������������������������������������$ H�dɒ	Y$�/��X

B��!F�H H������AАGdv�@��H����3&d̟���U��J>S��9NS��9A�i��1� �3���� t���� ,�e��f	���*؁�1�9NS��>�$�7�*�z7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y/fc��? dd�Ӕ�9NSdd��^# L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C7 �6�D'��������_�|T	���r��)�r��)�r��)�r��)�r��)�r��)�r��)�r���:�0�bbbT��R1I ��'����������$P(����9NS�d���>$*�S�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�e e�8X�9NS��*s�&G� �L�F�L�04
`h��)��S@��L�04
`h��)��S@��L�04
`hB4
y#�D#@��F\�����S? ��/�``�g>#L��r��)�r��)�r��`�]21���R*D�����dɔJ%Y��I$��	�&$H@�?��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�Q(���H�@�:	�/����000a&�p�� d�D�Q'�&L�d�G�D�@@!@�P}>�A H2D|��)�r��)�r��0Y�	�LҦ#�U#�V��nb� ,�e��̕@2��S��L�9NS��> fi�ȕ1T�ѹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��S��f��3�fr��)�l���+�b� �b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���P6�D'����&x3��Q�2fi�r��)�r��)�r��)�r��)�r��)�r��)�r��`� �����C(؛b
�?�����������dɔ
����σ��9NS&F��ٙ���Lsѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��) #/�2�)�r��)S��2< z`hB4
!��04
`h��)��S@��L�04
`h��)��S@��L���F�H�)��+�O�&g� g�8	3�)# 1N2O���9NS��9NS��*��#�H��!��k5�	���� �e���k5��$����2d�����������������������������������������������������������������������������������������������������������������������������������������$�2c�D�k5��@��������� H�B0*EH��8G��6"�@��/�`�"J%��P(�Dɓ��Y��lM��111��<�3LӔ�9NS��9NS�T#�08� :eK�y%���� ��X� �p�ɜ�)�r�����7�*�z7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y/fc��? dd�Ӕ�9NR4'�^#6�s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1��r���@&B!<dE\��g
�3�LT 3��9NS��9NS��9NS��9NS��9NR���">d��<2�Tʑ�8G��/F�Y��2������������D�����r��)�r�24����*�S�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�@��p��r��)�F p  ����S�B4
!04
`h��)��S@��L�04
`h��)��S@��D#@��S�
`h�eL|�DD3� 3�*��*s$F���:r��)�r��)�r���4΄�0L �&� ��
�R*A�!�?����D�I #Y��_±$�$�dɄ	���������������������������������������������������������������������������������������������������������������������������������������	$H@�$ɓ(�J&�Y�BA$�'����I$d�z*EH��I���P(B�U
���P(T��R
�ɓ&
��R*FTʙP
D,9NS��9NS����tS��L,X�,X�,zn3 `�dr��)�T 34�dK٘�&nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��T�(�� l��ٜ�)�r�#&f���� �b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���L����/"*�\��'��	�0�> g)�r��)�r��)�r��)�r���X,&	�a���ĩ"�)
B�$�'��������������"J���*��r��)�#K؂l��UJ�9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4�@��p��r��)�e$dfP�u�{��04
`h��)��S@��L�04
`hB4
!��H�Q�)��SP!�1�m3(`73�fT�L&/�(<�3�)�r��)�r��)��ʹW#%�/��/�blM�:��A �'������/��XBA��k$�@D�A�L�0�"x@�?��������������������������������������������������������������������������������������������������������������������������������������@�$ɓ(�J&�Y��k5�I /���ɓ&b�"�d�z(�J$vG`�d�zAАa&�H� P($O��$H���a�r8G���~*�\����:r��)�r��)��!N2> ����y�r��)�T 34�dK٘�&nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ �ə�)�r���ə�d3�g�@�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b������3���L�f �O���p��#&f���9NS��9NS��9NPygEAPga!�����C(؛b�� ``` H��������������$0�9��	A���r��)�#K؂l��UJ�9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4��\��c��9NS��H�̠!��)��y#�L�04
`h��)��S@��L�04
y#�O$x)�#��٨ʘ����"�*�����X&��σ��:r��)�r��)�r����3�('���e��d�z5��fY �$O�����H$`�:@�P�+ĒH�H2ɓ&$O��������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�H2�%���k5��c����	Y�2�̙�2a&� �:�xd�z
�U
�@�PQ(�I�&$O����(�J&@���2�P�f��i�r��)�r��)�r��)�r��)P| ��q�*b��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���@�? dg��9NS��34���������1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C73����"�D+�b8/f�ə�)�r��)�r��)�f��4f�S*eH�#��@��k5�&O���������������D��2�Tʄ����9NS�ɑ���L���	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�) #/�2�A�9NS��# 83(b:�`��F�D#@��Q�)��S@��L�04
!<�৒<���/c.L��E�&~^�������'�<�3�)�r��)�r��)���02�Tʑ�8G�A��k&L�������2d�%�(
AА_±$�$�dɄ	���������������������������������������������������������������������������������������������������������������������������������������	��&L� �e�J%Y��k5��?���&L�(
2@�blL��/B�U
�;#�D	0�SblM���"�f�Y��b�P(�f��"��L�0t	�U
�0���x�*��9NS��9NS��9NS��	A���n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ ����r��)�aW71##��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��+�$<�b����2;/"*�H���a�r��)�r���� �00�T��R1Q(�I�'�����������������1?��Py�r��)�	@1ٙ�qSG=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ�����9NS��9L��������/b�Q�(�hB4
!��04
`h�G��H�R:�`����B	���AL�A #>)�I�r��)�r��)�r��(<�2D|�  	�� @̙�2P(
%�@�?������ H����P(!F �:
%����2dɓ&$O'��������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�I�f�Y��001����$�/�a@�PGdv��؛�	056&�؂!�P(��! ^���$�LK��V'����$!HR3&d̟���
D,9NS��9NS��9NS��*��n2%LU"�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ ����r��)�2fiW71##��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0^DU�f�@��)�r��(�c(e�������������������$Ha�s*eL�P| �S��9@a( �32n �h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�A�p�
pX��9NS��H�̠!��F�L�F�L�F�D#@��S�
`h�eL��C2�� �3	�1~	A�i�9NS��9NS��9NPygB`�&q�LLJ�R*B��)��������&L���k�!HB�f�YD�Q&L�2d�������������������������������������������������������������������������������������������������������������������������������������������D�&L```�I�f�t	�D H�����@�$�A�I ���V(
d̙�T*�Pa�r�@�(

��6&ĩ"�b```�H2��/���D�
����X�`�&	��i�9NS��9NS��9NR����)
^ Џ!���y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���f0I��� 6FL�9NS��6FL�*��$bds01s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1WBHy73�"�D���r��)�r��i�@� ��D�����������������$0�9��	A���r��(% �ffM�M�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�2�0�E8,�S��9NS)# 0C2��#����04
`hB4
!��5S м
���rlʜ�Ɋq�|��:r��)�r��)�r����3�0���$	��6&��k5�&L H��������$����!HR�!HBA|_
ĒH�H2ɓ&$H@�?���������������������������������������������������������������������������������������������������������������������������������������D�&L�H2�$���kAА_±2d������dɊB��lM��6&�ؙ ^�ə3$vG`�lM��3&d̙�2fCC��f��@�P(	$�@�?��"B���2b�|_blLLL@�<3L�4�> g)�r��)�r��)	���? 0��A���ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ �ə�)�r��hN�\�ČL�f �!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���ON��r��)��`�3&d``c�����������������$0�9�2�T%�)�r��>l�8_�|*�S�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4e�a��pX��:r��)�e$dfP�u�{<�৒<�G��#��٨ʘS"�
g�@�����H�S����9NS��9NS��9BPy���0������}>��I����k&L�@�?���������,�k5�B��bB�f�YD�Q&L�2d����������������������������������������������������������������������������������������������������������������������������������������@�!D�&L```�I�f�P(k5���/������A�Q(�A�t$
�2fLɱ6&�؛bdC.��@�3�Y��
��R*FD2�˦@��HR��/��@�t	ɓ��d�@(
 B� ( �X,�9J��#L�J>S��*�	��,_�=	!T�٘�& �����s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<J�@E0� ��3��9NSdd�ҮnbF&G3 s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1�`D'��'���9NS�%��9�6&� H������������������ H�HR� �#��9NPJ����	U*��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѢ �z�69NS��9L���̢/2�j2�<�৒<���/b��"��� 3����� F|S����9NS��9NS��9A�i�3L�4f��#*eL���2�P(����2��������@�#�Y�0�8a�qHR�@�Q|_
ĒH�H2ɓ&$H@�!D����������������������������������������������������������������������������������������������������������������������������������������	L�2A �$�@E�|+�@�P(+
��2d������ɓ&k5���@I���"�T��eїE�AD�Q	0�R�T���6&���*�P�AА$I|_
�@�� d�$���I$���#�p�?�P
 L�2BCbŋ8�i�f��)�r�#86a8�B��=2�^ Џ�R���(��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���f0I��� 6Fpl�S��9M��3Ex�@ �L�f �!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���ON��r��(J> H2@�	������������������P(@� X,r��)�	@1ٙ���Lsѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�і	�B)�`lr��)�r���%s96g�4/�C*`E
�D@A3= �3 �p ����t�9NS��9NS��9J��d��� @a `�H�"�@�I ������������&L�D�Q�A�!���)
@�P(�k5�J%���dɄ	$O����������������������������������������������������������������������������������������������������������������������������������������D�&L�2c�DB@(
AА000$O������@�%�DB00#�;B;#�D1P(
�R*A&`j_±@�P*EH�
B��H$a�!ʑR*B�@�``c��$�Q(��8G��O��;#�D3&d́�xr��)�r����p�78@e� �bT�9���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��^��	1�~ �ə�)�r���ə�\�ČL�f �!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!��I&�`!<dA8/g)�r��A�?��@���"������������������"A@�Q`�Y�r��(% ��~	���Lsѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�і	�B)�`lT 3��9NS��H���و�@��ɳD'��%9NS��9NS��9NS��r�FK,bbb@�3�HR�?��������L�1����D��� 0�9@�P1)
B�(
AАQ(�I$� �e�&L H�����������������������������������������������������������������������������������������������������������������������������������������@�!D�fY ```�I�f�P(!F�Y��2�������&L�/�aB0(
H�"�T��(
$�@B�@�U
�T�� �/�c d���"�@�I$$O��ɓ&I$��%�$�&L��``eL��3L�4�9NS��9O�x���	�,_��!>T�R/F�E�7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���P3� ���9NS��#Bp�*��$bds0��(b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���ON��r��)P| � H2@�	������������������	
� ��S��9@a(�O�	U/��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ,�S����9NS��9NQN2O�����4΃��:r��)�r��)�r���X,Ca	@��blA�t$	X@�?��������@�#�D
�(
�@0�8�)
@�P(�k5�±|I$��	�&$H@�!D������������������������������������������������������������������������������������������������������������������������������������������&L�������|_
��:!HR�#Y��001�������&L���k2@� ^���V�#T*�P�P((�J%�@�g��؛@�P(
f�X@�?����I$fLə�4�> g)�r��)�T 3dd�Мe!@O/ hG��@E � ��y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y/fc��? dg��9NS��34W�����`b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���L���p���)�r���:	@��2� H��������������������@��`���9NQ�6B/�>l%T�㞍�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9��qSL� ��g ��)�r��)�r��)�r��)�r��(J>APg P
 O�����}
�|+&O���������ɓ$�@F�Y�R�"�@�P(
�@�P1!��H5��b��_&L H��"B������������������������������������������������������������������������������������������������������������������������������������������	ɓ&e�d�����D�k5��@�Pa�qHR�f�Y$�'�������dɒI "HI$���AR*EHB�@�QR*EHe��fLə*EH�!�0�8������� H���&&!0L����9NS��9NR������*�2�g# A�ĩss����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M���f0I��� 6FL�9NS��6FL�*��$bds01s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1WBHy7 �	�"	��{9NS��9O���2� H������������������ H�P(@� X,r��)�3��A*�i��J��=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���&�̙24���)�r��)�r��)�r��)�r�����3Lњ3@���2�d̙��@�Q(�I�'���������dɒ@@ t	��)�(
�@�P(��@�Q��k/��X�Q(�	Y2dɓ&$O'����������������������������������������������������������������������������������������������������������������������������������������$O$�2d�A�000Q(�Mf�X�!�1
���V$��"�������ɓ�# d�@�PB�U�2fLə3%H�#blM�a�sY��L�?�2dɓ&$O��L�1@�P_��_�x��`���9NS��9NS�2A���f����l��p�6�nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��%N "��~ ����r��)�2fh�������1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C7 �	�"	��{9NS��*���~2@�	������������������P(@� X,r��)�3��A��6�_��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ��7E4e�a��1� ����)�r��)�r��)�r��(J>�2C�9���R*EH0�9$�'��������$```�/�`P(b�P(
��@�b0�8�)
@�P(BA��k(�J$�```�H2ɓ&L�0�"���������������������������������������������������������������������������������������������������������������������������������������� H��@�!D�&L�H2���VAА!�(
�!��t$J%d����������,�/�`��H�#blM��P(2@�
����@�$��P(�$��AD���ɓ�
�R*FTʙP
DJ>S��9NS��9M��3AeTD ��=	!T���E�C �&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�8��a� #86g)�r��hN��F F&G3 s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1�`D'��'���9NS�%������$O�����������������$H:��0���S��9F|�%\�6�	U/��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9�Рp2�0�A�9�|�')�r��)�r��)�r��(l�0���$	����T*�!HR'��������$```�/�`P(bP(
��@�P(C�B�(
AАk5��%�$$�@D�A�L�2dɓ&L H��"B�������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2��H�k5���H�C�
�@�bBA$�&L��������D�I !HR�@�P:��@�P(
?�ɓ1G�3&d̂�@��"��$H���@�P>�O��$	">d��i�9NS��9NS��6FL��LU�\e��M��F%H�"�ds����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y/fc��? dd�Ӕ�9NSdd�Үnb ��P9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0"�D���r��)�#L�$	F@���"�����������������k5��LLA4�|�9NS�g͐�)̀l%T�㞍�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ������	�B �32_���g͐�T 3��9L�4�2D|��`���9NS�Tp���~?��2���/F�Y��2��������&L�$�5��b��)
@�P(

�@�P1!F �P(�k5��f����  ������ �e�&L�2aD��������������������������������������������������������������������������������������������������������������������������������������������$�2dɓ$�@E�|+��H�#HR���P((
��)�f�A �'�������dɓ&L�I�	0�RI$�$� d�#�p̙�2b�$	�&$O��ɓ&_±�2迋����<3L�4�9NS��9NS��> `�pA3M�DA6O�1T�Ѱ��3s����y7<M��s����y7<M��s����y7<M��s����y7<M��s����y7<M��s���P3� ���9NS��6FL�*��$bds01s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1WFA07 �	�"	��{*��r��A�� H��$O������������������f�Y�
���9NS���d �s4�l%T�㞍�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"�T�d�� �z��'�8,�a(T 2����)�f��h$	FTʙP<�`�YP| ��i�A�@(�?���p��@�PQ(�I�&$O���������"I�&I$��f�X�)
E�@P(
��@�bR�!B0�F�Y��k5���I �	�,�2aD�	$O'��������������������������������������������������������������������������������������������������������������������������������������������2dɓ&H$c�D�/�cY��
�!HR1P(�A@�P�#�D�L�?�������@�$��k5�&O��"Mf�X�B�؛b
���V5��b��)�f�������dɂ�@�B!� @Ca��S��9NS��9M��3A���l���BHU"�A���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&��{3$�a� #86g)�r��hN��F F&G3 s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1��r��ON��r��(<�3��$	 ^����������������������k111A�r��)�3��A*�i�*�S�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9����L���yK���0�6 ���d ���9NS��9D0�������G�,X���@l$*EH�
�D�L�?�������� H�dɒ@@ t	�!���P(
�@�P(��# P(�� �k5���I$��$���� �e�&L�2aD�	����������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2dɓ$��E�|+�f�P(!F�!��@�P(
�!�f�Y$�&L��������D�&O�000(
P�@�P( H�A �AА(
��6%�@``c��� H�I$P(�#������$�σ��9NS��9NSdg�'HP�g�Q���A���nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<��1�Lٖ/�2fi�r��)�`��d9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0"�D���r��)�r�@�$d�z'������������������Y�����3LӔ�9NP���9� �U1�F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4�J��h0'M�� #8�T�@J|�)�r��)�r���X,�?��,�H5��f@��B!��� a�rI$$O��������$I �e�±|
�C�
�@�P(
�a�qHR�!�
��H5��b��_I !������A �&L�2d��$ H�$O���������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L```�IJ%����t$�@�HR�C�
@�PP(!HR5��d�A�$O��������HlM��#�;@P(I �!��P( ^��x*�P��# �"���@�%�D��_��_�l&H��#��9NS��9NS���p�7�2��`3�� Nnx<��&�ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�� t�d7<J��E�ٖ/�2fi�r��)�2fh��d9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�b�2	����ON��r��)P| � H2@�	������������������	k5��LLEAPg�)�r���8 Fq�P8
�h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ������	�B �323@0��t�*�P| �S��9NS��9A�i� @a3&d̒@@/��&L�@�?��������&L�����+��P(�P(
@�PP(
�a�qB0�# P(k5����V(�J%�D``````�H2ɓ&L�0�"B�'�����������������������������������������������������������������������������������������������������������������������������������������������@�!D�	$I2d��,```�IJ%����t$B��)
A�!��@�P(
 �P(�Q(�&L H�����������@�P6&�؆�
 �C<6&�ؙ ^��xT��R(
�H�/�b����/����2f�Y�U
�T@�  �APg�)�r��)�r��&̱�`��SH�!���y�e!���nx<��&�ɹ��nx<��&�ɹ��nx<��&��{3$͙b�#&f��)�r�#&f���@g�@�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���ON��r��(J> H2@�	������������������Y��bbb��S��9BS� #8��J��=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ�����p�����d� J���9NS��9NS��9L�2@l$p��Y��$O���������$�2c�Y�B�
��P((
�@0�8�)
B�`
��t$�f����%�$�$�@C�A�L�2dɄ	$H@�< H��"���������������������������������������������������������������������������������������������������������������������������������������������'�$H@�$ɓ&L�2d�	$�|_
ƳY�

B��b�P(
��@�bBA$�&L���������I�@�B06&�ؙ�2fE�A�2��8T��R(
�@������P(J%d���� H������D2�˧�����r2#L��r��)�r��)�2fh,���� ^ Џ8�� T2���nx<��&�ɹ��nx<��&�ɹ��nx<��&��SH�2��6FL�9NS��6FL��1 �a �L�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���&BxȂp8^�S��9NPH���/AD�������������������Q(���f��)�r��)� �b�=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F��"��� ��S� S���g͐�|��> g)�r��)�r��(<�3L�4��
�T*�f�X@�?���������D�&L�I��H1P(�A@�P(
�!�!HR�# P(k5��f�Y|_
��D�I	Y �e�&L�2aD�	$O������������������������������������������������������������������������������������������������������������������������������������������������� H�$H@�$ɓ&L� �e�I "�D�_±��k�B��)�(
�@��P(�5��d�A�$O�������ɓ$���vG`�*�P�3&d̙ˣ.�blBL$���g�@��@�PlM��6&�؊B��H$���D�J%@�P2�P� @a3L�4�9NS��9NS��#A4�LU�d��F �<�R��ɹ��nx<��&�ɹ��nx<��&�ɹ��nx<�1T�ѳ,_�dd�Ӕ�9NSdd��^#6�s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�tdp0	��2 ����9NR���@�$d�z'������������������e��f��i�r��(J|�g�	U/��G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�@�U2�#%�$|��1�P� �P| �S��9NS��9NPygL�2@l&&&"�U
�HR�����������@�$�A�Q(�A@�Pa�r�@�(
�A@�P1)
B�(
�F�Y��k5�J%I$000000H$dɓ&L�2d��'�	�@�?���������������������������������������������������������������������������������������������������������������������������������������������������$�2dɓ$����I$_±��k�B�`)
B�@�P(
�@�P(B�D�Q$�������� �e���H(
�U
�T*�Q�6&�؛blM��5��e�|+blH�#�@��H����2d��t$
�T*��3��`�X,�9NS��9NS��> `�pA3M�DA6O��8|�!���y7<M��s����y7<M��s����y*b��fX������r��)�`��d9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0"�D���r��)��πH���/AD���������������������2��4�9NS��	O�pS� (z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���h�G=9����Le�a��&�̌�P�x	O�p�> g)�r��)�r��(<�3�\���H��������@�P������������@�#�|+B�a�q@�P(

�@�P(
��)�@�P(k5����V(�J%�D```�H2ɓ&e�d�dɓ&L�2aD�	$O'��������������������������������������������������������������������������������������������������������������������������������������������������� H��"B�&L�2dɓ&H$d�H�Q(���k5���t$
B��b�P(
�@�bBA$�&L��������```

B��(
��6!&`jQ(�K��V#�;C2fL�a�rA ������,�H1dC.��?��0���4Μ�)�r��)�r� �*�#0�  )V�	{3$�T2���nx<��&�ɹ��nx<��%LU"�l���34�9NS��34��&x L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C3�������p���)�r�����# d�@�?�����������������(�J#(e�4�3NS��9BS���6�_��F�z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѣ���hP8
�/�>3@2di{>
��r��)�r��)�r����3�('����}>�blMf�Y2d���������ɓ&I$����V�#�@�(
�A@�P(
�!�!HR�# P(k5����V(�J$�H```�H2��,�2dɓ$ H�$O������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�H2��,�H2�$�D�Q5��f�Y�

B��P(
��P((
��)�f�����"������$�I��H
�؛�@�lM��*EH�
A ���&L�I "d�����J%@�P2�P�q̑2A(<�9NS��9NS��6Fpl�qSaWpl��x�J�'7<M��s����y7<M���*�z6e��l���r��)�l���+�b 	����+� �b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���` ��P"�D���r��)�T 0H���/AD�������������������Q(���2��4�9NS��	O�pf
�`(z4sѣ���h�G=9���F�z4sѣ���h�G=9���F�z4sѦ�����p�����0�*��r��)�r��)��σ4�3Fh�?���p���	05(�J$ɓ���������@�$ɓ$�@F�Y�R�"�@�(
�A@�P(
�!�!HR�# P(k5����V(�J#�A�L�2dɓ&L H��"x@�?��������������������������������������������������������������������������������������������������������������������������������������������������������"B�$�2dɓ&L����$�(�J&�Y�B@�!
B��b�P(
�@�!F�D�H2�������@�"��_B�a�s dљ3&d�}>���!D�Q��@@ ��@��@�P�� �H2���ɓ&k5�͉�6 `� �0X,r��)�r��)�T 24A�4�d@��3H��F%H��&�ɹ��nx<�1T�ѳ,_�dd�Ӕ�9NSdd��^# L�(�1]�s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�13��D'��'���9NS�F��H���/_�������������������De��d���9NS��	O�pf
�T�d�����h�G=9���F�z4sѣ���h�G=9���F�z4sѦ���9/)����
s`�b4�*�A�9NS��9NS��9J��d����4ʙS*T��R1I$���'����������"I�&Q(�A�t$�(
�@�P(
�@�bR� P(�� �k5���Q(�I$���� �e�&L�2aD�	$O�D��������������������������������������������������������������������������������������������������������������������������������������������������������@�?�	L�2dɓ&L�H2�	$�|_
ƳY�
B�a�r�@�P(
�a�pP(I ��'�������"A�t$ ^���/F@���T��R*EH0�8@�?�	X�P(*EH���!�6&�؛bb�I��񁁁HR��R*FTʙQ!�0J>S��9NS��9O�x���	�,_�=	!T�٘�& �����s�䩊�^��b�#&f��)�r�#&f���A��@&C��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�`	��!<d@�f A�i�9NS�F��H���/AD�������������������Q(���2��2G)�r��)��P
����sѣ���h�G=9���F�z4sѣ���h�G=9����Lf�s=2B���P�x	O�p�> g)�r��)�r��(J>�2C�9���!�!HR$��Dɓ���������@�$�A�Q(�A@�Pa�r�@�(

�@�P(
�!�!HR�@�:f�Y|_
��D�I	Y2dɓ&$I2d��'�����������������������������������������������������������������������������������������������������������������������������������������������������������"x@�!D�&L�2d�A�000I$��%�|_
��:@�P�)
A�!���P((
�!�f�X���������$�a�sblM���"
�T*�C�I /��AАlM��6&�؃��HAА*�P�#�;@t	�A�L�0�"��$I$
����#$G̑�r��)�r��)�l��ل�)
��9xB<T�( EP�4�&i�ȟ �r��)�l���+�b� �b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���L���p���)�r���:	@��2� H�������������������J%���Uʹ9NS��	O�pf
�T�d�����h�G=9���F�z4sѣ���h�G= �R���L2ٙ�f2@ N�Д�S��9NS��9NS��> e\���ŋ����6&�؈F���������D��f�B01P(�A@�P(
�!�!HR�# P(�� �k5���I �$���� �e�&L�2aD�	���D�����������������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"I�&e�d�A �$�@E�|+�f�t	�`)
B�a�r�@�(

��!��H$aD�����$�P(bB�?�D�B���"
�dɓ&L�P(blL��/B�@��P(�@�������dɚ�f�blM�����⠨3�S��9NS��9J��F�h8f���Wpl=	!T���*�%A�9NS��6FL��1 �a �L�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���&BxȂp8^�S��9J��	@��2� H�������������������I "8G�W*�d�9NS��*��  ���yG=9���F�z4sѣ���h�G=n �hP8
2�2�8_�|ٌ� 	@3�/�)�r��)�r��)���0?���(e� d�:��d�����������&L�I�f�B0(
�@�P(
�@�bR� P(
�f�Y|_
��D�II !���A �&L�2dɓ&$H@�!D�������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2dɓ$�@D��/�cY��
�!�0�9@�P(
�@�0�8:��I$L�?�����D�	�� H�Y��lM��6&�ؚ�f��D��� $�LJ�R*@�C<#�;CblM��)
Dɓ����ɓ�Fd̙����@(���g)�r��)�r��A���N2����"l���r��)�r�#&f���@g�@�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b���ON��r��(J> H2@�	������������������HG�*�\���)�r�A~��*r2^Q�F�z4sѣ���h�G=n �iS���Hx/�>_���g͐�T 3��9NS��9NS�%�i�f�`?���#��@��Q(�&O���������D�&L��f�HR���P(
�@�P(��@�P:��Y��_±$$�@C�A�L�2dɄ	L�0�"'���������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�H2�	$�D�Q/��X�k5��@�HR��@�P
�@0�9��k'�������H$b��)blM��6"�@�0�9��"�� :��Y��lM��2@�J%�����$�@A�!ϧ��$	FH�� �|�)�r��)�r���9NS��9NSdd��^# L�(�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C7 �	�"	��{9NS��*�$	F@���"�����������������000G�*�\���)�r�A~��9/(�G=9���F�z4*�S*r2^QG� ����)���9NS��9NS����t��$��yə3!�!�$�2d���������$I2d�  :����@�P(
��@�b0�8�)
@�P(�k5��f��D�I �$���� �e�&L�2dɓ&L�@�!D�	�����������������������������������������������������������������������������������������������������������������������������������������������������������������$ H��"I�&L�2A �$�@E�D�k5���H�#HR�C�
@�PP(!��/�bA ���������	Y��k�@�Pa�r;#�D2@�&L�$��/F�؛Y��$O�����2f�Y���_��_�x��i�r��)�r��)�r��)�r��)�2fh�� &b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���L���p���)�r���:	@��2� H�������������������O�ҮU���r��)�T�f2@S���z4sѦ���%T�c4���f
�d���� �P| �S��9NS��9NP�|">d�sT*�P�)
D�H H����������	H$e�D
�
�@�P(
 ��!�!�
��H5��e�D�	Y �e�&L�2dɓ$ H��@�?������������������������������������������������������������������������������������������������������������������������������������������������������������������$�2dɓ$�@D��/�`t	 �P(B001P(�A@�P1
�%�2d��������ɓ&L���k2@�blA@�Pa�pB!� ^�  �����L�0P(T��R2�TʀP
 A`�Y�r��)�r��)�r��)�l���+�b 	����9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�f�`!<dA8/g)�r��A�� H��$O�������������������#�\�����9NS�/��d��	�=�A���O�1� �^ς���)�r��)�r��A�	A��L��$	����6&�؂�@�������������dɒI #Y��
�C��@�PP(
�a�qHR�# P(k5����V(�J$�H``````�H2ɓ&$H@�!D��"������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	$I2dɓ&H$d�A�I$��%�|_
ƳY�
B�a�r�@�P(
�a�sY��I$���'�������&L��)
F�؛blM���"�� �!	������000P(�����~	�`�F�Ӕ�9NS��9NS��9O�x��`_�<�ϓs1���9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��nf9@D'��'���9NS�%� �$	 ^�����������������������#�p��r2r��)�|��3�x��2�2�8_�|�3�% ς���)�r��)�r��(�*� �����C(��k5�ɓ'����������"I�&I$��f�X�!
�@�P(
�a�qHR�!�
��H5��e�|+J%������A �&L�2dɓ&$H@�!D�	�������������������������������������������������������������������������������������������������������������������������������������������������������������������� H�$H@�$ɓ&L�2d�	$�D�Q5��`�:!�R� ���@P(
HR�%� �e�	������� �e���H(
�@�0�9D�Q&L�������$�Q(� ^����� M��3LӔ�9NS��9NS��9Fp� "	���F&G3 ��r��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b����2 ����9NR���@�$d�z������������������$�8G� ��> g)�r��ɑ��ٌ� 3�e��૕��9NS��9NS��*��f������8G�P((�J$ɓ���������@�$ɓ$�@@�:C�
@�PP(
�a�qHR�!�
��H5��e�|+J%I$000H$dɓ&L�2d��'�	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	L�2dəfY ``````�I��k5���t$B�a�r�@�P(
�a�pP(I$���'�������@�$ɓ$�Y���� ``c�������L�0t	�U
� `��S��9NS��9NS�2Fp� %T� �^�&G`	���c�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���(���p���)�r�����~? ^�������������������������}	�`��9NS��*��T����)�r��)�r���4Ι">d��< @�R*EH�P(I "d���������� H�A �(�J �P(0�8�P(
�@�P(��# P(�� �k5���Q(�I$�$�$�,�$&L�2aD�	$O�������������������������������������������������������������������������������������������������������������������������������������������������������������������������$�2d�A�H$c�D�/�`t	 �P(R� ���@�P(
 ��Y�``` H�������� �e�&O��������$�1dC.��~?��W# �X,�">d��W#&i�f��)�r� �6bf���Ȋ�^gɹ���C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1]	!���r��ON��r��)P| ����2� H���������������������H/��/�4�3NS��9NS��9NS��9NS����t��$8㘘���T*�!HR$�@AD��������� H����Y��)
B�@�P(
�@��P(
 �␤)�@�t	�Y��/�b�D�I$��	�,�2dɓ&L�@�!D�	��������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�2d�A�000I$��aX�5��`�:@�P�)
A�!��@�P(1!F�|+	X@�?����������������	Q(�L��/Dp��0� ������C(�b��X,�9NS��6FL�¼ ���@�O��s1��c�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s���&BxȂp8^�S��9BPy�	@��2� H�������������������I
�T*��da]��t�9NS��9NS��9NS��	A�����!�2�Q�6&�
���������&L�I�f�HR��@�P
�@��P(��!H
��H5��e�|+J%���������dɓ&L�2dɓ$ H�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������$I2dɓ&L�2A �(�J%�|+�f�P(!F�!���P(
�!��t$J%d�����������������ɓ&Q(�D!�R�"���#�2�Q�#�H�9NS��9NSdd���z+�U*�3����3��s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1s�1�`D'��'���9NS��> `�$	 ^�������������������,�HAАGdv�����3LӔ�9NS��9NS��9NPX,@(�?���(e�blM���k&L�����������&L�D�QAА)
B�@�P
�@�P(
 �␤)�@�t	�Y��/�bI$I$��	�,�2dɓ&L�@�!D��"���������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�H2�	$�D�Q/��XB@(
�# ���@P(
 ���:������������������	��H$blGpygNS��9NS��	A��,و$^ ؼ����	�ٸ��!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���&�`!<dA8/g)�r���4Ο��� d�@�?�����������������@�blM��C(�b�i�f��)�r�����9NS��	A���f��4f�S*eH�#��@��Q(�&O���������D�&L�Q(���H1P(�@�P((
�@0�8�!�@�t	�Y��/�bI$000000e�d�dɓ&L�2aD�	���D�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�$ɓ&L��e�	�,```�I��k5���t$�@�HR��@�P
�@B���V$��"�������������������H3񟍀@(�	A���r��)�r��)�!8/`�{2�!<dDbds0��(b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���L���p���)�r���~? ^�����������������@�#����"��� 	��">d�`�Y�r��(<��C�x@(���`�4΂�`�$G̐��FTʙR�T��a�rHL�?�������� H��"F
%�(
1(
�@�P((
�@0�8�)
@�P(BA��k/��X�I	Y2dɓ&$H@�!D��"���������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��@�!D�	L�2dɓ&L�H2�	$�|_
ƳY�
B�a�r�@�(

�@�P�D�H�2����������������L�0��(e�<�APg�)�r��)�r���34g
�U��FX�0���s1���9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�f�`!<dA8/g)�r��A�� H��$O���������������"I  @�P3&d̐ @��$G̐<�3�)�r��)�#�H���U
�TdC.��?���A H/��/�T*�P�``I ������������$```�k5�B�a�r�@�(

�@�P1)
B��``
��t$�f����%���� �e�	Y2dɓ&$H@�!D�	��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�$H@�$ɓ&L� �e�I !XV/���VAА
�!HR1P(�A@�P1�� ``` H��������@�$ɓ$�@D�H�2aD�������L�0P(T��R @� ���)�r��)�r���f L�xa�EZ/`#�p0	��C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C�1�C7 �	�"	��{9NS��	A��$	F@���"�������������D�J%@�PG�?���4f�">d�S��9NS����t M�؛bI �%�@�P6&�؄�I���``001����������"I�&I$��f�X�)
E�@P(
�@�Pb0�8�)
@�P(BA��k/��X�/�bI$000000H$dɓ&L�@�!D�	�@�?����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	L�2dəfY �H2�	$�D�Q5��`�:!�R�"�@�P(�A@�P�!HV��A �'�������I  P(b0�8(
(�J$ɓ��������I "�@�G�?��\����|�)�r��)�r� �����*^DU���>M��(b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!�b�!���&�`!<dA8/g)�r��A�?��@���"�������������H$��H6&�،��2���� ���)�r��)�r��Cc?���Y��$O���������@�$�A�Q(�A�t$�(
�@�P(
 �␤)�@�t	�Y��k5���Q(�I$���� �e�	Y2d��$ H��"B������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�$ɓ&L� �e�I "���f�X(
�# ���@�P(
��@�
�%� �e������D�@@!��$�LL��/F@�� d�@�P5��d�H�2�������	Q(�L��/E�_�� �&�d���9NS��9NS��9M��3Fp� %\��e�� L�(73�9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�f�`!<dA8/g)�r���4Ο��� d�@�?�����������$�@B����"��$	A0L �fȨ> g)�r��)�r���X,�Qbbb(
	�'����������@�$�A�Q(�A@�Pa�r�@�(
�A@�P1)
B��)
@�:f�Y��k(�J$��I	Y2dɓ&$H@�!D��"x@�?�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	L�2dɓ&L�H2�$�D�Q/��XB@(
�!H0�9@�P(
�@0�9��k$��"����ɓ(�J"��)
��	05	0�P�	05	0�Q@�P(
!HR/��X``` H�������ɓ&k5����� ��`���9NS��9NS��	�0���UJ���dv ��P9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0"�D���r��)�#L���~2@�	�����������ɓ$�@B��)"�T��3���H�� X,r��)�r��)�r���� �@����8G�a�rd������������"F��V�#�@�P(�@�P((
�!�!HR�# t	�Y��k5�@@"I$I$��	�&L�2dɄ	$H@�!D��"������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��"I�&L�2A �$�@E�D�k5���H�#HR�C�
�@�P(@�QD�Q$�d���$ H�dɒI #Y��)
B��P(
�@�P(
@�P(
�@�P((
 �P(�Q(�&O�������000)
B��3&d�?�r�FJ��r��)�r��)�T 0Y�&H��xW���73�9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��9�c��n0"�D���T 3��9NPH���/AD����������L�2HP(�eїL��2�4f�">d��i�9NS��9NS��	A���*� ̩�2�D2�ˢ�@��Q(�&O����������2d�H�k5�B��P(
��P((
�@0�8�)
@�P(BA��k�b��Q(�I !������dɓ&L�2aD�	$H@�!D��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'��"B�&L�2d��,``````�I��k5��@�P�!�1P(
�a�pP(k5��%�$$�@C��/�`t	��)�(
�@0�8a�qHR�!HR�!H0�8a�r�@�(

�a�pt	�H H���������$��B�@��}>�,X�3LӔ�9NS��9NS��34'��/fTD'��3��s�1s�1s�1s�1s�1s�1s�1s�1WFA07 �	�"	��{9NS��*�$	F@���"��������ɓ&k5�́�/G����?�`*
�8�9NS��9NS��*��f��x� @�"�P(
%�@�?���������ɓ(�J �:!HR(
�@�P(
�@�bR� P(�� �k5��f��D�I$��	�&L�2dɄ	$H@�?�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�$ɓ&L�2d��,```�II "���f�X(
�# ���@�P(
�@�bR�!HR�!�R�!HR�C�
�@�b0�8�)
B�`
��t$��H�@�P(B001b�P(
�@�P)
B���k'�������dɚ�f�;#�D111��<Tq�r��)�r��)�3�L_�E*�Xq�2�,3��s�1s�1s�1s�1s�1s�1s�1s���(���p���)�r�����# d�@�?������������``lM��C(e���!�0l�S��9NS��9NP�|�0L8㘘��"�T�C����������	H$e�|+��H1P(�A@�P(
�!�!HR�# P(�� �k5�±|Q(�I  ������2dɓ&L�0�"x@�?������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	$H@�$ɓ&L�������$�(�J%�|+��H�B�`)
B�a�r�@�P(
��P(
�@�P(
 �␤)
B��
��t$�f������V/��X�/�cY���� 
B��)
E�@P(
��@�!F�D�H2����������2b���3&d�?�P
 A`�Y�r��)�r��)P| �f�@�"���dE\��L��?�1s�1s�1s�1s�1s�1s�1�`D'��'���9NS��� H��$O������� H�I$)
B��B������s$G̑P| �S��9NS��9NPX,Uʹ,X�����B�
	X@�?��������&L�����+��P(0�8�P(
�@�P(��!H
��H5��f�Y�V��I$I$��	�,�2�ɓ&L�@�!D�	����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$I2dɓ&H$d�A�000I$��%���kAА
�@�P�!
B��b0�8a�p��!�!HR�# P(�� �k5���Q(�I$�������$�$�@E�D�/�`t	 �P(R� ���@�P(
����:	$�2d����������I
���X�c$G̐J>S��9NS��9J������*"�DF&G3 �`s�1s�1s�1s�1s�1WFA07 �	�"	��{9NS��*�$	F@���"������2d�  a�r�T�� �<3L�4%�)�r��)�r��(, �@����2�Q�2�/�bA ����������&L����|_
��`P(�A@�P(
�@0�8�!�@�t	�Y��/�b�D�I$��	�,�2dɓ&L�2d��� H��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��"B�&L�2dɓ&H$c�H�Q(���k5���t$�@�P(!F���!�@�t	 �:f�Y|_
Đ�I&L�H2��,``````�IJ%Y���� B�!HR(
�@P(
HR�f�Y �e�	�������@�"��_ ^�������4�3NS��9NS��9NSdd�ќ+�	W71���g�A����C�1�C�1�C�1�C�1�C7 �	�"	��{9NS��	A��$	F@���"������"I�&Q(�E�A#�p�?�`f��h<�3�)�r��)�r��(<�A�@(�?���p��@�P_±2d���������$I2d�$���k1P(�@�P((
�!�C�B��
��t$�f����%�$�$�dɓ&L�2dɓ$ H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ H��"I�&L�2A �$����I$Q(�J%�|_
ƳY��k5��f�Y��k5����V(�J$�H``````�H2ɓ&L�2dɓ&L�2dɓ$��������D�_±��k�B��)�(
�@P(
 P(_±2d����������2`�P(�"�@�  �`�Y�r��)�r��)P| �|T	����	���^�&G`	����9�c��9�c��9�c��9�f�`!<dA8/g)�r��($	F@���"�����&L�k5�blFP�G��� �0X,r��)�r��)�r���3Lњ3@� fLə(
�D�2��������$�2e�DB@a�q@�P(
�A@�P(
�!�!�
��H5��e�|+J%I$000H$dɓ&L�2dɓ&$H@�< H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ H��"B�&L�2dɓ&L�2A �$�������HI �$�$�$�@D�H```�H2ɓ&L�2dɓ&L H��"B�$ H�dɓ&L�2c�H�Q(����� 

B��b�P(
�@�P(@�Q$&L��������```�P(�8G���L�(<�9NS��9NS��>�$l�8^̩xW##��nf9@s�1��r��!�b�!���L���p���)�r���# d�@�?���񁁁��U
�T_��_��$	r�FA`�Y�r��)�r��)�r�">d��@�3�R*EH0�9$'���������D�	YD�QAАbP(�I���P((
�@R�!B0�@�:f�YD�Q$�@C�A�H$dɓ&L�@�!D�	$O�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�$H@�!D�&L�2dɓ2̲A �e�	Y �e�	Y �e�	Y �e�	Y2d��$ H��"x@�?�	$I2dɓ&L�2A �$�@E�D�/�cY��
�!�0�9@�P
�@0�8:������"������$� ^��g�`  	��">d�S��9NS��9NSdd�ќ+�	W71c(�����`��Lb�!�b�!���L���p���)�r�����# d�@�?���D�J%��H�#6$G̐J>S��9NS��9NPX,Uʹ,X�����B�B00���������$```�/�`P(bP(
�@�PP(C���!H
�f�Y��Q(�I$���� �e�fY �2dɓ&L�@�!D�$O��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O$ H�dɓ&L�2dɓ&L�2dɓ&L�2dɓ&L H��"x@�?��@�!D�	L�2dɓ&L�H2�	$�D�Q5��`�:@�P�)
A�!��@�P(
��|_
ĂA�$O�������ɓ5��b�U
� `*
�8�9NS��9NS���P&/Ǣ��R�9{ ��&��P�1�C3�������p���)�r�����# d���ɓ&Q(�J��3&dʙS*�`�f���4Μ�)�r��)�r���:��0�ŋ/��/�blM���k2̲@@�?��������@�$ɓ5��b��)
@�P(

�@�P1)
B�(
�@�:��V(�J$�H```�H2��,�2dɓ$ H��"x@�?�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	��'�$H@�?�����"B�$�2d�A�H$c�H�/�cY���� 
�(
�@��P(��D��2aD�������e�	���3&d�?�r�FA�i�9NS��9NS��>�$l��#���p<�ϓs1��� ��P"�D���r��)�r�@�$d�z'�ɓ&k5�́�/C(e����@(�A��σ��9NS��9NS��a!������}
�Y��H2���������ɓ&I ��t$�(
�@��P(
 ��!�!HR�# t	�Y��k5�J%I$000H$fY�H&L�2dɓ&$H@�?�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�@�< H�$O'������$ H��"I�&L�2A �$�I$I$����V5��`�P(B�C�
�@�P(C���H'��������"J%��P(>�O��2D|���9NS��9NS��34'�쫛����d ��P^DU�p8^�S��9A�i�� H��$O�Y �
�������� H �@��`���9NS��9NS��A�3Fh�2�T��8(
f�Y2d���������$I �e�J%P(b�P(
�@�PP(C�B��!F �P(BA��k/��X�Q(�I "I$H$dɓ&L�2d��'�	������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�?��������"B�$�2dɓ$����I$Q(�Mf�X:��P()
B�a�q@�P(

��)
F�Y�``` H�������ɓ&k5�͉�6&&& x����9NS��9NS��9F|T	�p� %T� �^DU�x�@ g�@��9NS��> `x�"�T�  ����)
@�C</��/�#WB`�&	A���r��)�r��)�r�">d��H fLə(
� H����������&L```�/�`P(P(
��P((
�@0�8�)
@�P(
�f����%�$$�@Cɓ&L�2d��$ H��"x@�?����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O�D�	L�2dɒ	X���$/��X�k5���H�A�!���P(
�@B�
%�2d����������2b���3&dʙS*@(���g)�r��)�r��A��p`��Y� �4Μ�)�r��H��#*eL�R*EH̙�2@� <��4�	A���r��)�r��)���`�& @a111*EH�
B��000$O��������$I2d��,�k5��@��@�(
�@�P((
�!�!HR�# t	�Y��/�b�D�I$��$����2dɓ&L�2dɄ	$H@�!D��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2dɓ$�@E�D�/�cY���� R� ��!��@�P(1�� �&O��������"F
���},X��#�HF�Ӕ�9NS��9NS��9NS��9NS��3L�
D��Tp<�3�)�r��)�r��(,	�`�q�/��/�blM�:��,�H'���������ɓ$�@F�Y�R�"�@�(
�A@�P(
�!�!HR�# t	�Y��/�b�D�I$��	�,�2dɓ&L�@�!D�	������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$ H�dɓ&L�2d�A�H$d�H�/�cY��k5��@�P�)
A�!���P((
�!�f�X���@�?�������&LV/�� dщ���⠨3�S��9NS��9NS��9NS��9NS��9NS��9NS��9A`�X���~?��2���/F�Y�``` H��������� H�dɒ@@ t	�!���P(
�@0�8a�qB0�@�:f�Y|_
��D�I	Y �e�&L�2aD�	$O'����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2dɓ$�A �(�J%�|+�f�P(!�(
�@�P(
HR���V&L�@�?�������&L
!�� �X,r��)�r��)�r��)�r��)�r��)�r��)���0?���p��@�Pk5�ɓ'����������"I�,�Q(��@����@P(
��@�b0�8�)
@�P(BA��k/��X�Q(�I "A �$�dɓ&L H��"B��D�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$H@�$ɓ$����I$Q(�K��V5��`�:!HR1P(�@�P(1
�  2d���������@��8?�ʹW# �4Μ�)�r��)�r��)�r��)�r��)�r��i���y�#��@�Q(�	����������"F��V�A�!���P((
�!�C�B��
��t$�f�Y��Q(�J%�$�$�dɓ&L�2aD�	���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$I2dɓ&H$c�H�Q(��f�Y��
�!HR1P(�@�P(1k5��$�2d���������D��g�? q�2D|��)�r��)�r��)�r��)�r���:d��� @a @��3&d0�8���@�?��������&L�$�5��b��@�P
�@��P(�1!�@�t	�Y��/�b���$������� �e�&L�2dɓ$ H�$O�D�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�	L�2dɓ&L�H2�	$�D�Q5��`�:!�R�"�@�P(�A@�P�!H�/�bA �'�������dɚ�f�T*�Q 0 �9NS��9NS��9NS����a0L  	������T*�@�P���@�?��������@�$ɓ$�@@�:!HR(
�@�P(
�@�)
B��!��H5��e�|+��I$��$������� �e�&L�2aD�	$O'�	���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$H@�!D�&L�2fY�H(�J%�|+�f�P(!F�!���P(
�@
J%dɄ	�����������)
Fd̙����Uʹ��g)�r��)�r���X,&	�bŋ����6&�؃��H'��������$�2��HB@a�r�@�(
�A@�P1bB�@�P:�����%�$�$�dɓ&L�2aD�	$O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	L�2dəfY ```�IJ%����t$�@�HR�C�
�@�P(
�:�����d��������$I$�
����b�H��"����)�r��`�
D	��>�O�@��Y��L�?���������	000_°(
(
�@P(
��@�bR�!B0AАk5����V(�J$�H�H2�	�,�2dɓ&L�2d���D��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2d�A�I$��$�|_
ƳY�
B��)
E�@�P(
��@�)
B���k'��������"Mf�Y�6&������$G̐,3L�4 �3���G�
�|_&O���������ɓ5��b�`P(
��P((
�@0�8�)
@�P(BA��k5��e�|+I !���A �&L�2dɓ&$H@�?�$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"I�&L�2dɒ	X���$�(�J%�|+�f�P(!F��)
�@�(

��!��L�0�"������&L��``T��R1112�Tʘ����2fJ�$�'���������ɓ$�@F�Y�R�"�@�(

�@�P(
��)B�(
AАk5��f�YD�Q$�@D�A�H$dɓ&L�2d��$ H��"x@�?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H��"B�&L�2d��,```�IJ%���f�X(
�# ���@�P(
 ���:	$�2d�������$```�k5��@�Y��000$O��������$I2d�  ��k�!H�P(
��@�P(C�B��!F �P(BA��k/��X�Q(�I "A �$�dɓ&L�2aD�	$O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�&L�2dɓ$�@E�D�k5���H�#HR�C�
@�P(
C��f�����"�������D��������� H�dɔJ%P(P(
��P(
�@0�8�)
@�P(
�f����%�D�Q$�dɓ&L�2aD�	$H@�?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"B�&L�2d��,�H2�	$�D�Q5��`�:!�R�"�@�P(
�@�P�!H�Q(�	X@�?��������������&L������k�!H0�8�P(
�@��P(��!H
��H5��e�|+J%I$000000H$dɓ&L�2dɓ&$H@�?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	$H@�$ɓ&L� �e�I "���f�X(
�!H0�9@�P(
�@�0�8(
$��Dɓ��������������	L�2I$k5��!HR(
�@�$�LE�A@�P1!�@�t	�Y��/�bI$I$��	�,�2dɓ&L�2d��'�	$O���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"I�&L�2dɌI "�D�_±��k�#HR�C�
@�PP(C��f����d������������� H�dɒI #Y��b�P(
�@�PP(
�a�qB0�F�Y��k5�±|I$��	�,�2dɓ&L�@�!D�$O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"x@�$ɓ&L�2d��,```�IJ%Y���� B�!HR1P(�@�P(�!H�/�bA �'�����������"B�2̲A$��A�!���P(
�@�P(
B��!F �P(BA��k/��X�I	Y2dɓ&L�2dɄ	$O'������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ H�$H@�!D�&L�2d�A�000000Q(�K��V5��`�:!�0�9@�P(
�@�P(B�D�Q&L�����������$�H2���V�# ���@P(
�@�bR�!B0�@�:f�YD�Q$��C�A�L�2dɓ&L H��"B��D���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	$I2dɓ&e�d�A �(�J%�|+��H�B��)�(
�@��P(�AАI$������������"Ff�X(
(
�@P(
�@�bR�!B0�F�Y��k5�±|I �	�,�H2ɓ&L�2dɄ	$O'��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� H���&L�2dɓ&H$c��/�cY���� 

B��P(
��P(
��)�f�����"�����ɓ&I ��t$
B��P(
��P((
�!�C�B��
��t$�f����%�$�$�dɓ&L H��"B�$ H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ H��"I�&L�2dɒ	X���D�Q/��X�k5��@�B0�!H�P(
@�PP(@�QD�Q$��"����D�&L���H1P(�@�P((
�!�!HR�@�P(BA��k/��X�Q(�I !������A �&L�2d��$ H�$O������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�	L�2dɒ	X���$�(�J&�Y�B@(
�!H0�9@�P(
�@0�8(
(�J$�A�$H@�!D�	���D�&L```�Q(���H1(
�@�P((
�!�!HR�@�:f�Y��k(�J%�D�I	Y�e�	�&L�0�"B��D��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�< H��"B�&L�2d�	$�D�Q�b��k5��@�HR�C�
�@�P(C�B�:���D�I$��	$�$/��XB@�)
A�!��@�P(
�@0�8�)
@�P(BA��k/��X�Q(�I !������A �&L�2dɓ&$H@�< H��"B����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�< H�dɓ&L�2c�H�IJ%Y���� 

B��b0�9@�P(
�!�C���!HR�!HR�!HR1P(
��P((
�!�C�B��!F �P(�k5���Q(�I$���� �e�	Y2dɓ&$H@�!D�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'��"B�&L�2d��,```�I@@"�D�k5���t$�@�HR�!HR�!H0�8a�r�@�P(
�@�P(
�!�C��1)
B��``
��t$�f����$������� �e�&L�2dɓ$ H�$O'�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	$I2dɓ&H$c�H�J%���f�X:��t	 �P(B�!�B�#��R�!��B�@�P(
AАk5��f�Y|_
ĒH``````�2��A�L�2dɄ	��'��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@�!D�	$I2dɓ&L�1������I$Q(�J%�|_
ƳY��k5��f�Y��k5��f�Y��k5��f�Y��k5���_±D�Q$��D�H�H2��,�2dɓ&L�@�!D�	�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������D�	L�2dɓ&L�H2�	$�$�$��E�D�Q(�J%�D�I �%�$�$�@D�H```�H2��,�2dɓ&L�2d����	����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�	��$�2dɓ&L�2d��,�H2��,````````````�H2��,�H2��,�2dɓ&L�2dɓ&$H@�!D�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$O$ H�dɓ&L�2dɓ&L�2dɓ&L�2dɓ&L�2dɓ&L�2dɓ&$H@�!D�	�'���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�	$H@�!D�	$H@�!D�	$H@�!D�	�@�!D������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������